PK  ў,J               metadata.datS�(U�J�S04R0��25�26UpvQ0204�*�H�L�(�54�*	�L)� � PK[���2   3   PK  ў,J               0.i��e\����t���t7�ҹtJwJI�4*����RJw�t� �t�4Hww,��s��yqι���g��\s�\O�O� ����<�� H�xZ d Lttt4L,,Ll��8/^���"�#�"���"���e�b���@I�*���������EX\$�����"HXXX8/pH_�$�Qҁ��� �D�rP��d$����y�hH���$dT4tL,���d$dT44T��^��~ � ��:���(��� ]�Xkℑ��=�5	)93+;������������������������[;{O/o�O���|���JHLJN��#5-/����������������������60895=�;;7�om}csk{gw�����������?\H 
����#�32**
*����}�3� �����&��!=(�H�[���W���}�5#�?�����7��X������\� 
��� `�����_U�6Z�R�/\-��"�\fy��ˈ<[+�������q^( �B�Є+ǵ̆Y��u��<�	�^�9����P����_��+��R.��7qƄ�=�~���������Z���mGtZb{nK�C�����	����R)�h-A'��60��3������r�� �t�1F���Z�[͟�u���2S���@w,��&;�'�z�N���·n�K���Yd17���*���|п�
��ǯx�f��?qáɭ�Y�	J�9��.!֚_��9�񰧸���R��Ui���=a6R�0�$���i��ݫ���9��{���(��Q"}��|��m:�м%����D"�#����'��z��~�ٳd?���!�����������.a?Nf��՜�X�@S��f�!�����R���<�A�<�J��h>�瀞�|'w���� �]}.�'B8�G�7Ә���n"��ki:.*JZaN۫��q��}�l��W�xF���^DP�#����Ѻ>B9r�[RZ��f��"��QV�D����q�{h@285��hL;�C��8-s�<uâ� ��$����1�
_��/���K<wG��7{�P�Ht���.
�H���
1:����Hw���D@�7�9�i�C�p�z��dg>�TeVuu�Rz+�t��Tl�~���'n��P��f�6��K�4%���9���ȅ ;�wW���~��O���Ż��r8i�t_�o��u8EGV�nJ������U�B��S暙21�_f4��W������*�� ��*���Ȫ�����q��Ƣ�i����<\�3˷X`i�;۞�om<;����Ozr{���õoǣ!y-��d�'`�	���\TZ�C9�}����쿽�����_��:��"�1�$,tU��7�bTH�U=t�r��P�Ƥ�����jQ'�w�ai�i��3�cBf�.�o"P�[u�6"�n�� w����+�x���6�'�w�����4U_�R����5�=4ú��%=g!�rJ[P�ל,�F���Zz	X�����m�3 aǐ�Kݘ�k���>4�^w��k��=�,�<T�:��<&̹�-8B���k?�4^h�Oed�rUn�C�ÞT�x�d�A��Eg�C�j�=��O��T�&7��Ӣ�Ns���#���������_�ͥ��1���$$�'�����8�kh@���I>�7���C�������<3�����ۑP_��ʪW!�'S���J�+��w���K���\�_��b�[^S�"�����u����x�����[�� 7m�^�N��A(.r��Qۑ�<���ř��}�D9�"H��!��o�n5���^���j�q�?��+r�㿝��v�.Kq}ٖZT2�H˻u��� �R*շG+��پ�?3I]��Ɵ^��&̐aOb�oف �y��M0�����:~�N�t�^5�T��I1�=�Y��Dr��������5Ԋ�V��ƤZ}��G�L�L��.v7��2H7��#�1�4�Gc�Զ͛C�_a�{��Ni-�e9?�Z�=)$o��=������ԊG��'@�$ٯ҅�L\����� ����'`���3�Vkܦ�%���a�%%�6W�S�V�ɷқͱ���俷7���?崕�YE:/�f"с�e	�����l��"Z��A��,/Ѩv(����D�hI��{������Oa��Jg���S��4�i[�J��Uf��C(Bnt�5�+�$cj4?s��*"yKd��p%d��{� �_��k�����0h
5�FR �����Y���Ck-r����rM�E��l�O��7������B� ޡoC�2����O�?$4��vnOrh���M��N:wtISf?��Z�	Yt`��pK��;ae�id���v)c[Ly���w3o������:C܋��ʓ4Y��WP�M4��$e�O��]C�ס���7�	�+�X�����>�*�����rV�9��f� �[��Z�,OMv�n�:rY��̛JXY1ș�qqz���T���\Q����V�W2M5��vp+�m�D�W�Mb�>��)~AME��j�=�<5~�:t��]�խ�Ѐ`N���G���J`�a4"-=�W��S��h	ж�PЖ������Q����X�~)��$0���Q��-�V_ۨv��!j9Z'��n���2P�Ũ��u͸m3�࡞�gGz�R�����3���b�J&'֏)%�)`�vi��
iQC�����ε�6����K��;���*�M�2�܄O�w�}hV����],ϝ^[�ZS�cc����~�[c��ꗇ9aLΛA�W[?)|
U��
aJַ�в�^u�"���C�yq1<�Vҕ+'���J�=�Н�WfL�3]I�g�4J���U2�4_p�B��z���{���I��3PJc��ȫ�>���Zz��J�נ��*�ȴ؅6*�t�Z�3�m �t��H��������ǜ �m��ێL��F>�jڸ��!�v!%�m�L���V���h�lQ��՚g���M=�n0�ףW�1;(3�|�/>�%:���̞�W�3�r�F��CY�5o�8oڼ�����Z�����v݁�:1�:k�&Y�2:yr·��5��I3�&�����Fo�����7hܳ�J�<�"vf`�ͯ1����)�F�Q��^�ʸ9g$�Z輋=PSڪ46��C	ʚF/���.��e�}���?�4�݀;�E���蹾��yO�O�00Ū7��u�9��[�ao;������媞C�xؽc����cq��+0a{gUߐ�{x�O�ZX۟ejR���4�����n�>!:j���bB|?�唱b{h���	�J�66v�0N_z��FU�2Ǫ�y�F !ï%?�� Sð$�����~���f_��~�B��;��7HhZ5���O�<��L��.�)�-�N��.�z���z��B�=��X��T�qy�+��G�2�Q�l��M�*�T��.�(���`�u�}���𽁉絕������^gt�>A�ı�^�F�#zu=����9�;�0���n�#���b1�m�П-f���v��� ��tv�X�׶��
#vr��P���r:v�Y���+%�j�0�j�������dT�MS9��Y�\ t�>Y�O]�*E�3�P��%@���*	��a�����%<�'^�/�q�_cdغ�O�� -�\b�p�
��R������ߩ����Yv�F��m�i{�+/+��V4H��E��Q��Ù�v	�1��[�'T�c�
�f6�p�?b�:r���aEKCnq�y�¥G4�zcĘ�2,`&��-1b��o�	��e�� �6��|�J�Q����dj@�Ibb�>_���=��.�&��Գl��ڻ�#�S��J�1!� �慕�6��C	�s�-���4IҴ��%M����ki5p%�-�`���Dz@�W�'�xAS��&[�;��b���8V�iOM�T�d�>�@�8:d�]�.Tb��ӹ�&��q��>���1Ϝ������A��)i1�����	2��XnjQ��O�!�qvм���Žo��I����P��{B�ZY�����y�����/�����px�><�	�鿃k*�h�.#�KJ/|�-�`�4�$0_3z>�.�勧�xAG�j�j5�r
&��v���9�NM��Ú���ީ=z�qԁ���i+DK��W`�]�V�[�,^�@��u���g�^��&	�.ԝJv�,l���lJ�ʡ:��+�98�I�պ�z�>}t��%�al�H���:�u1����D����=M�����8���]7j�G�G����R����Y�%��J�2Isrݮ�PdQ�F)'�b�)��

��� ��ǛF��4h&S�|������Qd��O��W�,�y���&������ڃqNM���+"��]����@�{��"~��r��"}Al��<\�͑�Ȑk)ue�,G�X�꼬n�tP��a�����	%��� ����{j���2�9&F�@��GW�g�oҌ������m�p��5���b�ϾQ!9�r�0<�d�;P9��ȄI��*	=:|�z5�X�k)�����P�}��h��}㊱���-�qY�=��x'��>�\Ɲg	��T1ͷIҟ�l�v2����97�{�F3� ҧ�kx�5)��Ain���ә�6�4�OU��S���֯"����+/t|7iՖ)�)�J��F&7�%?�i/��>�_����kI��:�h��@K��"�d7���	�+#T���k�٩.6���U�P��؞�ϝ�lSg�@���.�O��ҡ���W;����$E߅r>r��j����"l�꽇)������P2̷����x`��1�Y�-6���kd����$=���^Mc�K�
��X:�~ ��~0�X��0�z��X�[����jF�\���4���8ȥh�{��@1�xu,��$���7�f���>�����u>?!�}Oڨ��Ff�Z�#�i�4奓�J�R�u���ڞC//�G�Єnn����Yql7�%��x�_x�Eɵ8�aX��%�v31�G.q9G��;���طL��D&~Kq2w�&��}k�,�����.i�a,ۮ:�+�J���-Urʇm�
OySA���o��r���U_vwu��7W�z��ۏ$��U��S(����ػ+�%�@��J9�0�뿚?oS��Z�~6�C���6i��~#��K����b�a�f ��v\�]�&�8y~['7��烻�x���7zj�e�J2�5.�������<6��{
��'c��5j��]�}���O�0�������0FJ��5�;8�G�Û����J�ǂ�1��;��M�s���i�������kyIj�n�����_�?쭟���HW�>4����V�H�wL��$R*�^~D4x@y�s�����N�}S�Ig"��=p�T���
:}K�0��p�)������	��r1�7�A���׎{~��m��H:w��-�N����{��&���-��^-������-�ߕ��ˆQ�tT����i����ѹk��4���/ŭ-�-z�Ǿ|��sQ~�/1��#ZGS@�
�x���x�>�d����?W�� ��$����\��+5Z�r2�:��\>�ޫ�%���7�ې�vCH7�*�⢸��bSF�[xP�Dsoth^��Pʋ�C�CFݖ+�}?Y��I����!���D�Ӛ��η[�[KX� ��V^T�q���*�"���qJkŲqqkM/�R_��g��E���Fa!�O��AU!L��(�r0�>@�z��*����MU��)ȿLG��X1�_����&d��>��U�VT'q��Z"��35Q��^�*ﲹ�����U� |�MQ�z<��X���d�EdOO�09�sL��bZ^����@�JV�|6;��\�:0��<���fj�t��!p��yvr���aߤ#�j��0�6��&3��ӔU�}���<�z�z��$S9໗���(�������*�6y.���J��Y�~`�x�\��--U���R�VᮜV�}x�A[j�Br�%
�)�ڊ'��t����_��rxU�`���< 2�s̨�x��VD���8[���/}�g�~+��_�p�o�'�,�sJ'�ϰ˜���6cϺ�r�:�+q�LV���F�_9��jQ��Uλx3�0�ߺ[;8J��CC9�[
���$����A�1x�*���dT�m��
��g���6�A�V)�V�l�]�on�:F�Ȓ<�?�iN��9'Ư�8�����j�혔�K}���ͽm�k��_
�Nӡ��ͮ��o�z�B�pN�-���ag�uu��i7�>o��㤸ug�߲�R�YSG�j�L6Q��d�y�=>-a�A3��E�rcfd@ܸ�$�}���g8���x��ޱ�V��h]��#�Ĳe_3}��L��1��0�*�ϪQ�.�h���J�O3�%=q�E�$�����?^?ԗZk�$�_K�e/k�4�$�*>���e`�$����6�r���xx�R�C��m����F�Q.�v+<�vo�����ywJł�1�y�����S	������U��J�i+f0hp��(���j�%8�}R2���fp����L|��#�V�cyqr��O�9�N�x�d���;�t�Fn��(4<�����:�ƽ�$�X���U \L�GK�ۢ�j�3eףj���6?R��jPs]V�{i}��ְ�g�qǌ&��>�!k'.�0�UD�ԧl��P�⤐�>i b���U�y�54��a���K4�1S.�O�ϯU�$�\e��JA��$NӔ$� ��ŉ�U��xy攢 ��s�ZiI�S�y?�z�׾'P�J���%���������d����ѐ�g�~����L_���b%����h4�Q*N�'G�w�rS�=�]����
�*�Q��5!����h&�K�Ju;q/����ֶ���%qV_}�u�A��."�ʊԈ��ڭ9�~�毠5)�}���v�(|!$�����' ��ۆe|�K���,�7X}�L��i�\	J0���'���2����b����Q!�)�~}���=i'�߳A��'�ڜA?Ł���IuM� ���jc.�-��fq^�bŮ/0��)]X���<>������7R>��xB���,_��@>�A"���r���=�	�:z�	�S���kD1o��?�~v�8$�_��]0���Na��������vyP�ٖ�=��k�'ṀL6���ޣ��l��.<�Ks{�i;Gw�ԋGWVY�b��OGu��%vI;`�|�~�=q��`[�[�SY��FB8H�3�_Oa�Vƀ�Cԛͽo�r�f�u_�\]�c��o���s�мÆO�KP�
��	�ry���[��T��y�6;�J+�GX㚴/�iUrI�S��/:r�'��q���K�M!`�H��:�%*�fח,���d��¶��"���𥁷��[%N�sNHWA?Um�����3���0���W	Ʋ�U�P��\�1:�Trs3m��j+���S�[�<�*�8���vYO��A�N�u(J��Tut���[��������t&�nz��=N��S��[z�P�Ġf+���� �-�.^y�[��+�y^���op��o�T�¯e�f��kC�(�tG���� ��j
��9X<�Ȕ�8hm���"�7M;���a�9�܀��a-���1��e�xY����`��O�(��?U|�K�ó�\|?�p[ޘj`�S&+E���r7CW�3[WG]�U�q+^\�t�! �u����Y��U2�]h�m)&�:�w.f�ʢ{�@�_���@�8���z1��;h�աS��[k��`QAw���*�W1tSP3��i���	�۽��w��������
DU�O[\C�{Σ����.+��m�Us�z�s����~TR�I����1�]Ej57�f��r�� ������]9���?SBRI�B\�ǂ�Ks�S�zi�gsG�cک~�$=
Q�)�K����Ub�󭊅�T]"&�q�䜎r�b���Z��YL�#BDV~�8��y$�j���!�~ӆt�*Y�\R9�U��d}�$kyU��������#�s%�JvRE��t����hyR�@l�[���&yS	�q�µ�NWF��H��$z8�S�c[�xY��)�T�<~�+��F���~�H�4QC�]Vp��O����n���<ׯ@������B^�7׊f�tk�V�.���ň�`�Y�[0{�pV�kt��^�PA��
� ��,�yET}��Wgwx]Ay+ᗄ�{*n��?���nc�T���:�����Gt����y@W1�����W=�+u t��
��|�ك.R}P�<����yoJ������Ӿ�9n��˂?�{�B���7j=������g�_���!t�������7�T>nn@�F������'#m��K%�.<��1� ����P]}lj�YQJ�l�.I�?�2�Le��	L���f.���i��Z� X�֤*�\�B�W-f}���:��L8	�T�s~DB��c@�Hz~����'2B���k�S+�q_Y�J�-����O� ��ѩ|-��Ҍ��hU/"ᶆ/���cZ����;Mq�n�Le�5�i� PKM��"  �"  PK  ў,J               1.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��]�6�h,�b����^��:eBt���Ǔ��s�KG�����/>��!o���|.�i��X��:�GZ���{����N�'�|�pi,��$�a[�C�~�I^?Y��w��S��r����?���%���=�8o��Ĕ��'�B���/�U:��a�
HɤY[���E]K� 	|���7y�Ī�i��(����K����3�.��+���2'a����z>�vf����������g/��.l	t`Ń���n������;%�M�_��
�m������B��"�"������
�g.9�D���7['��JJ�t	[L(�L�-��o����?��U��3Mʚ��w:B������Nj���;eֵ�*�7v؈ �j���-fNZ�L��ʸ������俟Fq�/��V�����2���ʌ%3����<��u/���3L��.��[PW$�'�U$�q�X̜t��
�a��Y��[05N�M�]�`�DX�}Io����ʮK��x����=l�*���Ӥ'�ZJ]���40A1W����Wʫ��:���z��;E2�p˞B֜z�s�_��l���IH}��{�;���+��+{�3���g���ِ�A���l�.��\ܳh�쥰�?U�>�6:)��:�q�����翮�Ӌ���6)-4=���H�A-������l�W�09o������E����a�j�b�����~�_���&���G5ޙ�Jf�.ϥon����@���Z����6˙�r��ӸҴ`��#vI>�Y�0���ʶ|��|�yƢ�ԉ/nϺ�U�\X�לS��KZ��e��o��?����o=��,��������D�T/=ex�,����Y�\�5.��t���	 PK	r��  S  PK  ў,J               1.vec�UoQ�=�r��������Ci����������.A?�4�"���=|�sfND���'C�2�(K9�S!��hV�2U�JըN�$��f-jS��ԣ>h�d��٘&4%�fМ���lEk�Жv���lt2;Ӆ�t�;=�I/{z�}�K?�3���0Mb�^�\��2��3���I��}��1�e��D&1پ)zS�iLg3��l�07��<�//`!�X�����i6V譔W��5�e����4��6�[��6�����b�����>�s���0G8�w̝�Op�S��g9��4�B����%.s��\�:7����[z��;���y�C�X��S��y�K^�7����齗?�O|�_��ww�#���/~��'-�PK,�5�p  �  PK  ў,J               2.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��]�6�h,�b���J��b��<�����۱Q[��(<�����kb�g^��5S!�?�{��x����ſ��e]����/��^�`Q��|�FYs�덪��Ǜ_����q]��BڧU��nf/�p���nz�]^���b�&~$�-�M����?e;5W��<}���!��5�n��c$�X��s���/�����ԩ�T�f�x{�n���)��O�����ݖ��P�)~�S���H�c.�E��ٖ��͖31��}X��P	tx��㞙o6ߍ����T�mL��Wj�M�{?�o�����[7e�ɑsE]k�D]�ᬘ�%��J,c/Z��\-�[o�v����#��%ݾ����w��T�nد���x�ܵI��@_Ht	`ăY�5.�\?}R���!E�6s8}�o(����!jMܫ���_O����ɿ`����Qу>x,���n���1B������)p��#ua��IOZ���+�OIy��׷��Ʉ�i�'�*�������s�q��hΰ�dܷgr�)���4V���s��-ټ+rQ��>��g�3�SR�vVw��w�V��c`�BNj�ﰹ��b$��z�:Mz#�!G��hP��޹g��HK�ݔ��)ɐ�r[����yb�\�\���+�v�����O��?�r�IqP
�99��N����_��z>�/{�ӿ�$"�����N?<��}��`Ǵ�_����y�^���̊	k�x���=גw���U🎾qf��J���ϭ<�?jw��w���g��ړ���Tu�����\V�Ʋ���r��N��3�_�_�u�ᗵ+؎�>���߂k�mʙ�4J4����q�nj�ݖY%��8B�����7�ٮ���B]����	 PK')  H  PK  ў,J               2.vec�U�VQе�w?[�[�[������������A�Q*�!�����b�����W@�B��(�(�"J�%)Ei�P�r���NE���BU�Q��LQˬM�R��4�!����lBS�ќ���S.ژmiG{:БNt��=]�nt�=�Eo��7K�����d��P�1�o�)���(F3���c<�h�$����2���`&����b���������,a��2���
V��լa-�X��c��Fy���V�����ۥ�[��^�������8�]���8�	Nr�Ӝ�lq.��|��\�2W��5�g��F*���-ns����>x��Ⱦ������%�x��轕��|����W��[d����W��PK(�l  �  PK  ў,J               3.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��]�6�h,�b������8�Cn�z��޳͘'��?p�q}�K���ٚœ�W럪�n�ѳc�����������h�).�E����!#ᥧ�>�;�������1ˏ4ξ��?Û�{��i��d����|��Ϣ�Eئ�۝r��ū�uޖU��b-�U���	�j~���g���_i���%��=�E�xs��/�U�>w�ϓ�ϰ6���d�	_���lm���n�*���fk�_}�x0��m���7W��ԯ��Ƿ��0ε�
��JJ��P�5���7���w:R���x�.��V�@V<XJ��gO�޿���l��蟛����g�tMtO΄����/km�����+��l�غ���+�Ek]E�`֗����e�X���ت��:�X�J���Ε��+���˵NiR��M�CޱM��K�LwMZR�}��xƢ.6�@W�Q<r��ݓ�O&9ȾN��;��祡۷�.]:�Ct������%=�6i���]_�F�uJ�y�ꈹn��Ƣ%ui0@1�ֵ���G#J��V�m����W���k�9�����1�]�y!MN���+�z>�đ4����ww����|iU���;�c��t��X��]HL�DH���nߦ�n�<I/�����Z{�5��2��np|����Mʗ���$<�7X���.���fz�ѼeL~����g��δ��ʝ���y���x9����]>�\<�����Z9/"����=��n=O�B���[/���y���E�^���<}�U��B��O�;��~]����8g�i��V���j���lŏ����n*�x4͜q�S�'y��Fnͽ&��g��5;��9<�Ԝ�eO��*�� PK��{  :  PK  ў,J               3.vec�U�VQ�u��>[�[�[������������A�Q�9�|���7;"���W@!9��8%(�E�2KS����<�H�,��*T�թAMjQۿ�u�G}АF4��NS��iAKZњ6��
��ٞt���BW�����AOzћ>����f1��ʃ��2��`�ި,�hyc�x&0�ILN1ž��4�3���b6s��
c��͗��E,f	KY��z+�U�fkY�z6�1�c��fy[��vv��]��ۣ�W��~p�C�G��{�Op�S��g9��q!��E����U�q��LEqK�|����>x�#�=�{*?�9/x�+^�)�wz��|����W��ݛ��?��o����PK�e$�l  �  PK  ў,J               4.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��]�6kh,�b����q�)����{a\�G.��b���_Z�K�v�릢�0y�����;~��عI��_�I���(�[ԥ�&�U$�f_^�y�Ɲۖ���R��zꏻ�Ͷ~�g8�]|�Җ�����mS�����Ǫ?:�'�+��T�f�i֬EW]K]E�a����G�<�r6+����GY���R7���ϰ�j<���go��ʋ�6�+5��������R��}�V�%�5�@���O�-�O���-���O�}m����l�y�9�w��G���Z}����Y����c�s]EW��:��bg�ߚ�΍Q.������"����^����[7�0�����I����>"ٞN���"�_ɬ�*� �ʀg�g%o�j�js�>4���5�H�2�P0s_����}���I���s=�T���^��*sŽʩ���6.$*�x�c��z8�-p���]����|%i���y���Z�Y�DtgA��>�סI�ﲁ�^9�K|�����^�_&W�E8�D��g�bL�!�nB��=����>��d~n�r���f�?^��7d���<�o�t��Qs4�'O�{���P��9�ɫ�OX\;��pr�9�g]��2qGC�d��Z�ʖ���F������z���w�gX��T=;��1}�+�?�=gީx}��_�{�k~��9�����E7�ꃲ�7���[�ު�9��ĩ��W�ڒ������5���_������bE޹�.�egY�'�.ia|b�򟡂��iT�1_���3����5����ޞ��|��_�Q�M�ɓְ��TZ�E''��!��r�Cs����-���� PK�|�C�  4  PK  ў,J               4.vec�U�a�g�P�ۃ�؊������q����Σ�N��G��K�����wf"�$�?���S����tQF���@E*Q�*I6��jT�5�Em
��d���G}АF4�	Mݧ�lNZҊִ�-��^v�#��L�ҍ���!{ҋ���/��π�IL��fC�pF0�Qv����c�x&0�ILfJ�����4}�>C�d���\�٘�~�,b1KX�2��"��J�U�jְ�u�g�lL��n����lc;;��.v��۫�c?8�!s��i�1�q\?�INq�3����.$���_�2W��5�s���︕��~����>x�#�=q�S�E<�ż���$�ؽ���|����W��[����W��PK�)V�n  �  PK  ў,J               5.i��ePL����J	R(�AZw--V�Z�%XqnE\�x�-E�w��4$o�w^�r?�{�;;�3����vw�gv�
�RWQS�� 8 � P		��@ 11	-9))�JZV&v6V&a>.An��R��"�����|2��O�	��?�wbbb2R2rr���,�O����P�( 
�p� ��8x�8� ��s��� �%\<|B 1	�߄&* ..>>��觿q >5�NQEBݷ@.Oڧ!I�D�Ju�������Y{��<�g`d�}���$.!)%-#��⥊*DM]������������������>�~�a�#"��c�SR��32���)*.)-+���ohl�������gϯ޾����ɩ�ٹ����ͭm�������������_. ����E���/��	�����u�o=i����*%�}'��;����C�G|���_��$����"��������}<<j p*���:�$�ƨ8��!�gl9��e�JǛU�1��d�!5��HT��&rCcV���^Q/|=��ҋ `�p��C0��V�P��[�� 9��ٓ�2a"��b;g��Tϯ������?�%d�n;����uX�L��V���Ȗ;��%�����}�d�t40�͹Buk����{f���)�c�m ����5}���7h�۰�P�ĉ]{��Os׭\q���vV�Nm�@�v탉�t�^���#�u�\P�r�J/�dԈ1H�2�����*�=�g��ԬZ�`�L�1�������p���:��a)��HG�d�SkP'�e*aIYDm^O�N��:`�J������PٶVɸ��s��X0Q6{���p�?�:�@��Dx��d�L|9a/���Veh�g��i�+�)�x� Hܭ}㤭k%�f}�8��k���} X%��949�6��8�f.�j�]��;���ǌp��+�s��Wx�ME���{h8sT3�!_�;r���N�-vΡb�R��l��E�|\�,h>�Aǿ�(�LL�9w�
`.��-r{��.��٩�K����0)?�b~���'�{{Q�F;�����E6D�s#*Ń��0p�t���$�k�G�f�XE��K"O��LW���?�B�%��ʳ���gf���&���}{��lm���L�ɹSٰ������ꟸ
�QizuO�3#�qgv�ؽ�)���N��M�v�����D��\'[{�r?�{^	�X�??��c'�J#8̒Yt���JH�����.y�����a�C[��D�\��X��)�j�F��"��^�[h a��6�׆%2җ�,�����N��y������Ǎq�C��/��AZ�D��"�ť���N�]�S�$mu��xu۳�� a�o��^Ym^�l?�yW��n�5��r�]�o�G�ĸr7&f8�_'Ǐr�] ~BR�wen�ޅ���c*�i��l�k�GS3��þ�3h	��;���QU��n"�����<=49^���-���Oo��]�RH}h��6�֍Ku�k���M��gG�-"����#ρ���oҳ^X�4��lAP%'y��i���ugn�6i�sS����(���Ny��ʎ1xl���w�}6��7�x�Mqp���}���{s���;!�1���/�>i��;AYY�����^x��r�#{-�	������!��zf�ީ9Wfu��pJ��"l��>�\��+�S�U�Y�'R ��Ln�8@'���1}��~��U9�.��I�;[�����F�MZ���0Ch��W��B�;����ฐ��(9I&�_�v�ͯ��xn5CGc<Y��	��.����Vj��޵x�S�MU�xѸjψkA�������(�-%�����ްµ�{�so��ԟ�ۊAs̞h�H�w*[~�ʤ2N�Ү�[NDK����Ť�/��i�x����o����(����X@��ZV�����\�G���*���UN}�� !��|�����j����0�D��_-��~���p�C�����%=�m}w�`�A��F	��oG]��Lݚ�%���e�W�L~�wm�I-�_8_�����2���i3��;H�l�c���F��82�C���ںݥ�1�;�c�Ҝ��$��M�9���#U/(�h���z$6�L�B>7����`��ۛ-J�k���g��^A�X3s��es�q|��eA��f� r{^m��&��iG(�\�'���fPhmg����#Y��������u�X��������)���!d����?{��;�Y~6ɶv/��'c�ړ�I������Y���� ��Ω��`Y|!�藆��]��k�/<���֊�g�U㌜�J^6��D���/lz�Fޯ��)%:�9ci򏟜#<:i/�b>�e	x8m֜e�&U(��/��r�Qe��1��͌v$9S�2�!ib���i�úa�:-��2Ͼ�,�~�rE����*/�䰧��B��D�����˽��d��������=J�Ǚ"���� ����D����n�cJ�O��􎻗=��s�A�����Ts�f�ֽ}=>����!�>2���j0���������O�(������zUܞA ����T��^b�l��-@r��3*v3����_�W{�]²����&�m�6�:5�8�s�?��\XB��,���F�!4#.��N����wp��Q�M�)�V�4�M�iV/ ��a�?Ee4��
zSk� ��ĩ��B�˞S[B1�S�!�:n��)�6�j�!�Uan��u��!PBN��Ct.g"��*FK�_��PU���RU�T.t������fzc����`O(AKމCX��.Sn���Xj9̡?�i]�����OB�Vl�#.]�V������Ыm��� ���a�d!'�#:{�1�蓑��L��������P����J�s�Z*�AH��@���|LS��TFdϓ��#�`�=���R��]YG����,������}pQU�yS���?J�4Th*n>�B]���i��^�v�[�պ�nkX���r~��c��2�,��ȭF��o�V�r?ao�Ԧ��?WC��yubkٗ�Z��u�>��u��X-'�뛚����S*Aog��]�[I7E�����_�֤.�]�L�$3W���uϫ�EZ���^�/IY˨��{��t�	1�*�Y�駁�I�OHN�ߚ<]qA._�+B4Ë60p����F�n@;T{ӹ�$����S3��E U���9Đ5�����A��TՀ1`�'xZ�ߵ�;�F���>������5J?C-R���夠�M���k:��r��5�� ՙ��4�k��(ɶ�W���l��=�ƍ�w����<���o����϶��ı	�!б6ou��5PCJdK&|[�4tzfh��Q4POﲸ��/ȑZBhns��Ή�K_�4&�\=vdJ�s�[���u�����po�+цJlE;��wI�ܐ�`�'f4=^d1�.��IR�* P�|С=��(I=x��Ø⻥����NjpH��ڰ�\��N�T �|���4V~�zi]���g�����a�F3ћT��D�T�A�2[]zPY.��ib��w��굉����6F��i������vk�U��;%���G��)T�7��o�n� ���o�O��t):RY���(�t�] �w��@~�Sy�h���F�� ~2Y���n��=h4�OE��KN��L�P��3J�k�'�2k=W0kX�*&U�Y�Ɖ$YeQ�|������+��s�i�i��+��N�m~	��Vs5m�G)��֪,���Q��n�
�3#Ti�[I����?��c��g����i��
�	��ѓrڦQ��
<<�Y�E�kQ�̔�ɩp:����o��\��p!ZO���J?�9n�H��S��\�5P�+nS�{h�iΛ�θ���㋳��Zc�����@�~��[ս��7ˌ��Tw�_Ur�F����M9_k9_I���/ґD~��_-���9i@q��z1x��%��Λ��U~��w�����@�=�]ȇ{�W��	��*��}�F�rQ�BO�Wm����np��7��R�\���=�f�l)u:pM���q����;��}m��)%U��)4- ����>��=\�`$�j94
=|���R�y7�$�[��o\y��N�r*�HI��Z����@8�*�5��/����za*��3l,Nj�O���Q*�[�?�����z@�FJ��%�M�.�F w�D`���tR�C_5ҧJ�I��ms'fX�7
�4�)�?���f��'���:G���u+���oI�#K�_�p��Q8��),�.]�����Io���(�f�C���_K[:���vEl��o ���~9�<�?�	���cv���䓘�=_�Jr�3�z�u|�k�^���c�1�\H#QU����5r���%�d������4�><O�O1N�<"��OK[J��c��o��f�,|����f�����){o�ƮI1�;?_�7Q��iz�$t��-�wP�㍣���:�Ћ�I|�r���@7E�H�A��1d��e5f"�	C��p�/�Osk��iiO�ؤ�G���2���s��G�����Y�f�C��c�zM>l�X��<�����o&
�G�F��&��/\s���<�� ��xn�#`�_��KKXx�=���J��/{1s��,��1�j?;}
�V��wh
y�-K�[-�,B�x�+�&��>��>�n��:;{o�m�'�ʲ�afå�n��-�7����(<�xݖ�;�g�Z�P�ʂ����\��~��3h�zOw�7�@+;�7�J�܆�!��$��M������1��B���F�%��T���&?	pqv#�~ԩ��621��#`��G_.�%���/m��i|޿@����o����MM=2�I/�DƑl������2�H�B�A�4��!�e�$J�� �+Ɣ%����'��]w�u�K�Mʩʭ���t���d��}�m�!���U����4�s�)��,��
O��G���q��a��b೎�Z�fʕIP�8��<w~r.Q�~���.j�د=��BSJ�b�!<L�Gꄭ�ভT���q�lM��v����o��6b�ertdR��Ob�LU�����Y�<�RQ�0@�b�7�JdrV{d�K3�O>Q ���7���q�[�]�<wc@q ����Q1Ԭ��d������r�E�f�w�%NcU@,Aq��ϜBF��E�CF\m��75
n�7��rm�&`3t��R?? `?���u�	Z��k��H�Y���Z�sR/� +%�1�����������i&�i{[ާX��
8�6��vH��Vkh��`z�-��9ܶC�):3��A�p_�߾E7����(Pp*1�X��N�ۇ�f��1��}�R/*���u�O��
`x�I��r��ph���p��{����������F*�\�=URHc���)|�ɝ��V̮�{����2l2P��*�ܲC��i��{�D<�7���j��L�2@��Sxr���j�J�Z���sI�b�������6<�0�D����d�d��T�tȅ<�Y������<�Lh����T�k�Ϡ
�l����b|�Ⱦ(㒤Q@�zo��$�z��qY>���G��TWk�����8���,p9J�@��X I���G��x?Ap��QL��@� ����,D�6yߺ�&�:�E�C�0v,	��Q_g,Gnh��6���`eV�����m�V����iLKt��?��#�3W�7��Ut���f3PFn�����o-������}�Qc���Ȏd��Wq�>���a��O��b'��TO���KR�I��������!���:��2�`�f���e7ʜ�`I��ML;�%�ܸnfd��ޞ~8�RWV���\�V-6�n��=�^ ��H���Է3�U�1����[�6�Z#��l1\m,ާ���Snox�߮��霚sQ}kL�� 氜��]~vT@:�=��A��<�P(��`��c�[zNa�8Zv�CL۬�Ă�y�ֽ��mT�]�nY�'�]�>�v������k���C� �9��mR��c����A��&��t���������~T�+1+�h�j���p OeЕR>���+������N (i@~�/}�< nZ&Pq<��Aoó{���
��S�B����<G�O-_	�P���L(>�4�1�íʵ� `DW������U�'�w��E�X|��ywrl	�I��	��*RN�I#l⾄���\i��^�{����*8�?k:�-�Ӂ�p�����'1��s���������!�*�,��P�Z�m�՞;E��D����~�D�l��s�G��7�_���h�?�w�V�ޓ���1V��y�-챐0}Q�����s7e��Nk��82�YC�*�$���%n̤}BL�Jy�?����]���,>�[, ^J��nU�%_Ǝ��t�9o���I�P��<U`��E�����1��{�����ԉ]��}/��=
�&ؗt���v�&����D���+e���5���>:��~��?xcn.4	�g����C����ƞi$���1U��Ob�#�P�i�Y����~��FL4�p�3@+h�����Anϊ�n�,����ՅҔ���4ƾݝ:~z��$<��ReO�G͠?�*��rV&��L(`�f���5��`ߠi�	KH=����ՏX�@��M�_��/���xTk�{A�z���/dK�\��=��w|jџ������:�B�)Nq�C���˛�1��f��y�Dg
�����6n����D���`8�v�4?��x��j��k�g����ϛ�P�j{N�_�ܚ8u��h)+*#�.~�:��B_x�X@� ���YR����2��	Z.��/t�LU_��630�Tj�����%�}�S)bC0ݳ�4gG\�Q��t
ڸ+���V�S?dk�--���1�ni�f�_�S�KI�&���%¸��2��RcJ敠~O�-�l߆�P�H�ق�;�"J�]N���?��kȸd��R���)^
C��Y�JaR���@9��C���^2'GnJ�5S�<�'�
ڣ��M&)����Q�@��6��)�*������M��R��ɧ�ɠs��un��6n�Vdn�o�j��/y�E�v�U�(�@� ݽ��J�r�GC>�V6gX j�t]�g΄�;h�w�%p�&����M:�^��f6����r�g3j�o�^�F�[J�l��E}縄�So+�ொ
�+�]Vy2^if�g �����>jVᴽ��ŭ�,l��H�Y3�I�R0���p�bڢ{S34������j�h����ۓv�Y�Z�ΰ�ޙM"��qxl�)�������>vm�eu�/J���C.�C���M-���mJ8�!���]��;=��Q�P{��3�RJj(Y�������O\ �L`.��2pm��7L��<��Z�\�ui2ߧ���n$�ƭ�+�F��x�?�1�a�ZX��vl˒��ilP�y��q��2�5d���sѴ�����rQ����X��5��gE���G�\�<k�,xx���S��)�)�)�ӧz�m��ɔ^V�3�N:�;�sb�AkW6Wᮨ'!�����kR���js�I�p�#m���I
�+�T��Yy
����t�6�=��9U6�Rݝf{	d����a3�ZR�Z%��� C��Ce�N+�	������u�'���~L�0-��r���M�l��;� ��F����y�����pu�%�  gtS@�Ι\�V4���n�l4���`�9��$K�r1j��ßP�~�,�4��+j}��M���C���9/�i�(����Q�S&� ����xG�6]q\f%����k׆�3v�^�#�a�:U�[ H�����T�W��
`C��������OVa�'7����"�QiL|�ֆ�=$2�WJ�{2����i�k��|�6f�c��� f�8���O?�-ovL�u�1B�>N�2��A^�Z�W��}�ӱO�+�%vy�!Es6wi>���!�Z욐h ���&}��z?��,�F��)j�ʒg�\@Ӳ!Q�`��f�"?Y����Ŝ�]
ܷ�OmKd��f�E�6�u)d5��PU������YO�ߞ��a$��D��!�h�n|�b�ݦ�e ѽ?��5KW�&�E� ճi���P1�`ą����Nn��^����}�����T�/Fuc�ʹ�c�[�=����)#�;VB��U��:%��A�K7Mh�/0���52��|�M�A����,8�;�Ɇ��u��Y�j�^�����	z�:�Xf�z0�|�����e~2���*F)���\#��b��?��<��#1�M�����G,2�{=R���ڿ0:T�/���#������3E�2a��w5��v]��O>�,.���gY��?*�5�ٹO�M�u�E�s>���@k9Մ�&�.Hj��?{n�	5���wUF1�l{\M�����KmMh0�z�#��[~O�ɧ萏��l�nc�Q[q����cE`��P�R7���>�h�%>s4����m�^�k����U��E���k�,,�@�2__�S'Q	����y��%}�����%W�Q|?��M���c�O�������To�PtE��"v�? PKrj��"  �"  PK  ў,J               6.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��]�6kh,�b����=]����,�	�l;�;�������������|��wOv��P�_(z��Cb�&�����cJJV&ʼ	�m��XԀ�j��K,���3���Կ�z��������>�gXpmy�s�k)u�k[�w(�g�:�����Ɇo��ߢ�vm-H�w	`	t��e�����lh����_�y�9���L�ϐ�j����6��6�8��I}��Ǔg�9�c���B�t�W�tkW��"���pު[w�`��g����q������A����?���������%�~������a�5�G��ui'
'Yы�$�jN\����o��������s��˶YLQvK_�g��
���ה]|�7�T���W���
�V�V0ui,��y�O<��{�����X�o��ܤco���_��ʂ��hP�:)�	g�.�7TWy~m�]����f��d�"��Q<���ꍶܾ�U����f/۞�͖�V�{b�&�"��s������z�TA��c�{���^/�����X�`��.(f3n}���}���SfN�������������潈ڰ��τI�{�[����5o��e+.|L)tV~35v	���Em���u�������9s�l�e{j��>����ޥ�J��E_K��a�3+�d��m��{S�u����4��~�����V���ٓ2g=�wn�^�ȍ�J�A��Uy.��i��*~����9���kW֊�g0x��º���������yꢫ�)~�<�;n�w��3���+�G�̥�Dz���in���6K��l�mw�{=2~���X���\���]�q[��'��h�Ξ�]3�U����M PK9➇�  ,  PK  ў,J               6.vec�Uoa�����!8���CqwwwwwwwwwrA�Q,�l��\LV#R^$��s�|
(FqJP2eQJ��e)Gy*P�J)�e�R��Ԡ&���Rԑu�G}АF4���i*�ќ���iC[�v�=�H':Ӆ�ts��=�Eo�З~�I�?���@1�!e�a7�7��fc�x&0�IY^LNS��Lc:3��,f3'��\�7O�����,a)˲�Xn�B_�*V����c=���h�I�������`'��v�������� �8̑,��8��'9�i�p�sv�SA\�/r��\�*׸΍�(n���os����>x�#��vO��<�9/x�+^�&K�����|����W��g�#�����Ί�PKI�x�m  �  PK  ў,J               7.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��]�6kh,�b����H���t���#�7*ǈ	=zt����K��L?w�1�|�{:���_�񟡓�������5ǔ��L�y*�̥���U>tY�����C�b��1����~��������oQ.�;�p�|��+����Ώ襁��T�f�YѬ��4�M d�U>����*_4>�_g���j~<wfN�$�!�n����rMo���/M>�n|�W������l�|��hâ.|��<�?�N�;�S�/-���̷�w����[��gC��G	�����>f���E������y?�0f��X�@(�+��>#�:Q8��ɣ�ٛ8/=xB���Uv�ӳ�6O�����?�וߍ8��2�p��KF�W��U	�����:��R�7X_˴AWd��-�S�'��M���3��ʃj�l\�%h2��r޸�U$H �U�a�b$�����[%�[dZ-�����ퟣ�U=�?�������*7ެ�R����I�������e�g��V���޸�����L�԰��tE?��^�k���ykf�J{v���5F�ӛ���s��
��}�����9kv��yu�M0��i��R�����ߞ���n�=������fk������w�UJ��?�l�üOf{7E,��H������ڶR�-��)�Sv޻!�ok�/�i`����-�4�L|��R�i'��������C�j��a�:R5/�~i؇'�6�J)l��Z|j�k��q��������t��J�7�ի�<�z2zʋE]���o PK�$j��  �  PK  ў,J               7.vec��nUA Й�^ @���Cp���ݭ����k)R����Q������s&�	!����咥�)C٘B9Y�<*P�JT�
Uc&T�թAMjQ�:ԥ^���l@Cј&4�����lI+Zӆ���=l:�Nt�]�Fw��ᬞ���C_�џ�à�7և0�ag#�h�1�`�>��L`"�����L�����f2���a.�r����"���,c9+X�r�*���
X����l`#�R6l�ۢoe���Nv��=v{����9�Aq�#�X
�x̆�INq�3���`w��~�+\�׹�Mn��p��~�{��yD!����Oy�s�y�K^�:�������|�#����z�o��{H�?��ߩ�PK�Xx�r  �  PK  ў,J               8.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��U�6�h,�b�������6?�>lk��j�;�	?2z����������o�z��i�y9����6�+T�_�x����)%����4�mj��X���8{ ���^יI+~�c��$�������ǳ�5�m��X�9�]ў�V�����=�?���YZW[��m��*����ʷ��V.1̟���?������w����`��M��>>g�>�ʶ�?Ú�~�b���v�g���]���x�.�@BH��d[�\*]�Z\q���������Jw�T?6�Y�b�|��~q�٦�3��g�u�&P� cQוDW� F|8/%����֠}w&G�:��6�W��/C���.��Wfaw;�?C�Q�@��	��X��f͘	�U��"x0c���-��ɽ�͂�Bw�G��X<������޵3�
j3���[X�\rLv��X�ץ�xDb6�'��+�>����=].�`����ia8����h���2J*�υ=���|�����׃н��eV�+%:�>6J�ԉ������Ż�/{��.�$�w���K[k���>�x:�����q�z���L��i��A!�?~��%K��|��g2r�f>9�o�������w�i�[+��q�0����}�>
k��

ݎ�jV)�<h�c?O;=�g�xS�C�;|�;����!80��"�>�۔�_�2$�L�����?Ѳ��/?��>:��[����گ�\z�,�Z+_���Ó�f�L�oWq\���e�"��m�خq�UTu��� PK���  �  PK  ў,J               8.vec�U�V1���f���Cp����������ݝ��e�f�쇝��6"�E���9�)�E)F�E	�$�(M�R��TpNE���BU�Q��L)j���C]�Q�4�Q�Ec�	MiFsZВV�vW�-�hO:҉�tqWW���AOzћ>����_���d��P�1\o�0R�h�0�q�g����"&�S��4�3���bv��9�o�<��,`!�X��f��Lo�����b5kX�:�g�Ao����la+���v����-�a/���r��YđTG�c�'9�i�pV�\ʏ��.r��\�*׸���ݔoq�;���y�C�Gz��'<��y�K^�:K�F����|�#����z�o��{d���wV�PK� qp  �  PK  ў,J               9.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��U�6�h,�b�����<�nr�^������\��(YX�����76ʊV!��y��ed�?��d����-r��3l��*�uc��E]�k,��`���/ژ[����T6�2>�Y��۬��A���3Ȯ��y�wu����o�����\5��z��_� [LBW��<}���D���x��,��K���ϝl-��m�|�xf�ޖ��u�6�vinھ#>���[�����l���!u�����ҭ]E�si,j��͗&�m���]�f���ʚ�yg���3��:�����<�w���Z��ө7�v����[�I�*�4Q���B�]R����������o"_o�d����w��cJ����{��&/?S7�X}̕[������X��s�ϺSt�L�,��4w�����N�gL���n���$>w�)�
'vU�v��*
�Q<��5���Qo�W�N�~KfG�"gϷ��*�x�-�.�l�Һ�ׅu�&'�rH�/Ⱥwk��sˏ99M0�I��=��5�u�Tbė�ϊ��O}�{h���ǓJ:ܵ��_���V?�yd�~�غ��/��E+U���>Ww�ۈ���[lO���kl0�k��<��i�wWٓw'�g��:���k��s*�3�'L����Ytk�Y������)���u[���pYі@Wc�ҝ�[�b�N,q��#S{��뮝Y�gr=ݳ���B^�_mk�+*�a[&U�y$LU��������ٌ�fѿG�?W�
���!?�>j�.G���E]����	 PK��ܥ  �  PK  ў,J               9.vec�UoA ���^ 8���C�R�ݽ��Kq������@�Q�f����sNv��b^�����d)Ei�P6�PN���De�P�j�S]֠&��M�R��1��!�hL�Ҍ洈��R��5mhK;�Ӂ���$;Ӆ�t�;=�I/g��}�K?�3�R��aP̅���2��`$�m7����1�	Ld���Ԕ�9w�>���b6s��<�LX`W�/d�Y�R���)?��[��fkY�z6��M)6�mѷ����`'����b���>�s���0G8�B8��~����4g(�,�R
��.���e�p�k\�F�n���os����>x�#��vO��<�9/x�+^��=��{�����g��ov���!����7R�PK�Vpp  �  PK  ў,J               10.i��eT����0��"�"���CHw�(H)!C�H��ݝ
���"-1�<��u��}q����{���g�����v������� ο`E��� L�O����I��HIHH(�ȩY!�,���l������9��=��*(""ᖐ�~,,"��Mp���HIH����0?��@A�#d�p�\
�����������	��D�$����8 .�_�ݿ8�G�O�@P��J��A-��C��;���1���{1-=#�C�G<�"�b��%$�+)�����ML�l^���;8�=<��}���������)9%5-=#'7/������������������Go�����ɩ�ٹ����ͭ��_{�'�g����o�Å�p����\��p��@x��p����'��� �����](��Z!�k�w"a�ck�qbZN�u�����7��X������\ )���( (p��X� �f�͸�V�i���F�>E��^�b'�M�9��x�I��YTQ.��Gq�(<%�~�C�b�����2%v/�X�QL�����yR��s�Ū̴��u�>b�^P�pg:�`��Z?��� 0F�XB�AU�L��$sSf�z6�G�_�X�]��U�fF��Ӊ���w-Js��+�X�9Ge�����Ǝ�!�t���,�k�!�լ���f��k��5��+KH �|��ӭ��N������VS��5'xB���bۼ���&��:触���֐^��X {6y޽������.j�|��['�?R��9���в��7%��B[��O������/Ho���8��g�Xuw��2����a��Y�f��_X`�e�H�=�-|�����*b�YCV�.�:?����G�{�}�X��v|ȼ��2U��*4�B��o˰m!a���U�n��<Ӑ���Յ��\:p��u�;u��I�g�ҩ�}h`�3�6J�ʇ;<T���>��=1ٜɪ�5��2�$cyn�Ra,{U��K�%uk��D������/�o�Y�QJЦ��y�o�:�l���=���ޟ	/��Lw��J�=�U�V��G�����[��5,����g�p[������i��1ߧ��T��j���8����d�����%Q�������g_���I1��C�:���Aʹ@��tt����E���/؈�ڥk�_�X��M��<m�z�M~I~�H ��3jW@��&b�c�X�	��,�����<ܒ��-�ҟ1���b�����6�IX��8��)qHA�?#�vk��*Ӱ�/�x�'���If�l��ts���yN<�i�o]������{���|���ժݫF�����Z���XS���	OPb��>�0S::��F��7�{eHw�1 jtwWѡW�(�g���w��_-Z���.�(�����|}kD��7�j�$�B��8wl�N"?<{� �i3��<eR�VZj4�@�y��w�+c&[����9�~�0�C�8k��c��.j-�5f�l��=���h�p�%^��=e|�"�;�)�]����~���5N+�`�J�[�1������������ny�����>Ts3��˵MD���FC	@�SIhGk��]J�y�ar�X�f�&�H����`�ú��k�w�Kf�'7-�~�������'�(lwl��|+�;�e�Ef��O��ܮ�	��B�'�xϳ񙃵e� ��06f�	� t��'7j�q׸
�-���n���\љuEߊ1�8�h�@ўG׼�0o����=m ޮ���T���Yo��G=6�[�Wk�^;-_:S�J���d���>
�Liyo��l3�	V��M��92���5���}"�#)�o_��B=01�#���2�݌?o�� �N���+���_�s"y�`��Ak�f+�����@���r&Y{R��ׅ�m�7�~C��;l�˘��j���;�bz��6p �
؊�Y�R��i�5��8�7�>�w	Mh�(�����a���х��*�M=&�5�\�^��>sT�څ��:9�gm&b8:�OT�y���H�D<q.{*=�/�)ݿW�gO�/�A\$�7�DVW�q7HP�L�G�\M§>�&8[${�4f��.A����c�@܏޻)�.��tARb�/��P���&�w&,0�������(o��S���bd�����^�I1?K!��@Ld85�����;�*=w��OS������e�ւ+�����~i2�BP�t���s��	�z�asL�߽�`��V���	j2IMOb�P��le8;aG�K��M�%�[�n2��}�����4$K�����mʎ�}_�S�Eꙙm�����K�/?�Oج7�[6�*�P+�2�k::�*q!?�~�5ˡ��8�W]�
z� �q�Pz:R��d>d��2� �r���Wc[�-(�-�>կ�%�[Xg�kF+|��I>�Č��%����{uLW�n��R�f`cv��W;Έ
4L;@���J:LYe�2��ߛYQWA���c���B��T��"���G�ͱ��	,����p9��m�n�c��v�L|�����W�!Z���N.�k����j\3�"K�1
��u��r���^%�f��b��2��):�4��:�iW�RB�nZ0�{]�K�m�SÜ��|6�5�ä9X�ⶨR���p��3��k	f�8i�rR���{޻�;	U�����T� *���<1KL 6EgWmM�R�-];�	X���u���*C��]i&�?;vG�Yx���Ϧ�>F�����8�%E�?��{�G*��}��T6uƝ3vv��}��K��9�)S�玮\��ѭ���Y{HHN��3u���,E���8�M̗�n�!��l!Pm|��Q�k��D�D_n��,|"1�g�SW6ڱ`�fk#	m��
 �nE����L�	��{{9ck4��BssQX�ADv۳���(�nn��ޓF�wo�/�v�TS��fJX���0�6�W�>�a�?���#�^?`��}'���c��4l/�g�´UB��%/q��/���O80�x��8������;�mlpF�ƶM�!�N�`��g��{[��q6�>�_��W~U��&���T�|��\h:P��8K�>o9<��%��N�����J�.��U
In�2��1�R�`	_a�v���֬�ڢm���fy��u�yܺE��_�L���Ω<�����#�f�ؒ\8j�s[�P����ۏ执���l���6�~�
�|;�̉��mά�!��T��WÏ�A!~��
T��q8�x^���1��v:E�4�#���U��إ0��<��\f��g�۬�ϳ���^%�Eʉ׼�&i������zQ�&2n���AŢj��ՠm>��ޱb��/[��y��Q����}ِ��4ʂ?��K.��Z������_𱍓�u[�o�^=��'�շ�T��ך�{-���Y^X 8�@�q�Q+'�Yک��M��w��R�u�i�[Uu5S$%i�/5�bT｝��gl������6��'cw�D6!��1S��QB����Lj���n�l�w!����R��+�=�.��Z��{i�L�O�h�3v5�l��報t�����ҥl1���dw��N���c�W��obG����HES�s��L�!�8�;t�(�����)��}y�;��]�
~��G�_�p���.0����M���������O�W*LW��4���7��G2HO�{�̲�J�s�bI�h�0&p�[O���ƚ�3�.vb��V٦)�I�W��d�@y�K,�ɯ���N|��Qy<��;�2.�y�v��I�_N�.�q��b�����i��5"�Pn�[����q�^�3C�X���W�kG�dq��.T@���C�96���HZYg+��f�b�@�P�³V�s����WD	)W�Ĳ�(Q�/�b�g�%7�S��'��۽�)��3���`����Cu�*�/��������*�,��B���YKU��O���
�]�T5h_l|�ʜ��%���,Kc�@�̊�.�$��#�����-�l��/�Pm����zU�����X��W5O���A��y�$�17�O�
6�#�"UGd���QM#���տ-����<C���m���sZ������pPѧPm�b�h	ݾ�	�z�Z�\�I@����%b��V���IH��~8�x��ۤsB���~�h�yը��Q�}?Z y롗p��¿�'.�g�6�0�s���Z�U�&������qm@����򎥊-S/�W�O��x�d�����ɛ��9��U�-�y޲m$)hKS�x���+4T����"����Ί�<��fIJ?R):}�
?����a�s�Eg�%�I�k��ZG�lK�"L���Y�c�[Ji{�N=%�:�fX��&Du�mb�<S�k�t�c��Œ/ ��SVޅbrxb�d�J��i��x�٢T�D�<T��l�Ϝg֡z���~�*;�Nj����.���k}ľ?�y�~�8�ٳ�蹏�q_ãI��S5h$4��3"`�CgÇU\�y,-c�pIp~�9ˀ�=��1hv�<��.I�]�ut����P�:�Ёf��~�B}�3��2���ޑ|��Z��C��/�w-�Yr`f�|��9�9'r�Pi�o	hn�}(�l�w^�����6%zi�gk�����[��7��"$
L0
sK�]���N��bk���$�GYpg��<
�q�sykmu�����ˬ���N�[�;r�6�e(�C}:����i�Ϋ�Ի}�`���Bn3'/4>/3�$�����Ю��q���-���M-�1�c�f��2�@ޗ�I��I��S�\7��p��k3���P~�7���΁f%,����-�ʈ8��Ma7��9�g�J��	����yCޏ@)��?N�^���K�ϐ�g�]����A{�냀ھt*?��=h���[mo3榳@����y(v�1�,b��L�c���̔:ǚ3�t��g�E��p��Ez�;����V���g/��q�`a\N���Σ�;C�ͷæ�Li,k�Z��DM%�`Dgl��3����<���^���şT̀63&!u�-�;x��\ƸCw�{�/���"���'#�+�eQ�e�e�CT�>
�ei�����f}d�麒��ܗJ���!:*ԩ?�����������Ρ�o�z%�Q��PL	�燡�V��([�OG�Q6o�4�G#T�b��<�`�ͩp�[��'de�E���LI���e����rҷF�*���r���=7o��,�>URi�(Ȭm����_�>�Ypu��t�{[c�lJ�l�Þ|砿���Ҕr+�����3S\�z?�&�f�S��L���6W*��d0��n4��:����K���2��5|v��JMp�~]%'@�m�Z��y��h�X>7��raY}P=�C��-�k�7f�,��<�ǃ�M��v0�BW�o�j�Y���-�L���mMç�$���m�I�e�l{��ȿ�RL�-�hrx��.�>^�[m8��o��J4`�5Ț73�BrG�9�"o��w�lt�ľ����}���H�#޾dF��H/^:�ﲩ��T��~�yR�ɨ�3�`�L�ݻW�ڧf�b������C�N�V��,�2>�Sq�]B6�7��>���O&�߲Z�G���y�{�4�oX[4G�1@uԳM<Yd��R��_y�F�?%#��tɋ+w���4k}��
"����m��9�-uv��c�^|�.+WЌ!!�FɎ��	'��9��zB{j�ʇz�Z��%*x���A�8g��7T��Q��ߑ]��#`6c&��=J�_�xי�f�[NEz���������!�&�j�bB�F�M?��7�}�����@��)��ݳ���b.X\�5I�J����L�[òW$mӐ���s�7�*�e�)�K�5)��һ{35+J��ag\i��'0'y6�tR��M^6�pN�mV�FF��ΥK[��Z��TgH�e���جv��*P�OO�����/Q#2�v=���*�x�,ΰ�4��B$�^z�=}�~����؇�;����O�H�S�V;X�!yvk�R��,
;�ȵ��|�xGg\R���O��/<	���:��)�����kE��KS�Q��U۝�jdkIz��=������5��ǂ��.���ؚ9��@"LdH�K�Eg��LTG����I$����'�~���9��1iD�{a���
��b��cM�D��/!�D킿�mo�_�"�J�e��,����R%��ç?���E��̪��=�)L�}����-O(�t:Tr���|�%9+S�,��\��#����0��n��U��`O�y9�wk�Y����B��т9du�T�ν����<O@���,����4R4J�g<�9	��ۻ���Z����NG!3)r�bﭨpb`2����$u���*�/���iP	(7lVk|�m���:�9Bu�Z��]NE��k��A�����RejE?y��z��O&�B��Ǖh�dT��c��k�,j���HïF�*���e�r�S�0��vm������Q�8�d(���W��ɖȅ~�ݿV'gl+�gu��ST�]�J�G=VO*%[!{O�h6;�������v��D�z�i�a�:�9��Yg5��T�%mt/m�������6��َ���ן��e�c���V�`;��ʘs9L����@x�c�	����U�뤗��b�&���l���G~����Gn���V����AV�OF�8�=�w��~\	�.#O2\���|��0I�ʋ�L� �"�Y^N3�d^LL`M�؏�~߹>�J+���}G9O�:\�d��ܤ��m^�.<WDG��|�O��Y�|�p�i`Twۼِ2�kh�|_8�&���Ax ^���I�M���6�h���5���X�ܬƺ{Be�b�����y��b�G��L3� ��1�8�#�,��F���d�:��U=��;��:U �Q�x1��f��3����X��=d�_��梘�=N������|%�|yA���
��9�=�v!䰧+/z���ﺐ������ϋ8���.�f��Azę�\3Q6��1�c�Q+�(d��|+>k�8zm�p�����˙�r��:�O���<�%��N�"�u��±�Ė"��f�s�b)�q�
��7g�п��J6;���h�*LN�C����2yX�[{�e�K��7]��	���$BԂ�L�����.b���;���˴��f��
�Ԍ�Zmêuw49����y���i�R�Դ�h�4R2��r���h����.�)|�x!����P���7�
fi(�/�yiȤ�/^�2����ܟhc��2��vewԯ�`T��S�����]�F2����~.ڜ�l�E�:n(��ˀ��χ�7�W��J��}n�T��^�6oaD��'�����2Ӑ�M���*�2��tTF&g�9lZe���si��ȡ��&!'�O�LKڎN�����l�3��F!w���%�y�ǂ�p�p�iM���?�@��c.e��^��;7ԁ����Doeo�T�����G�T��&���c�7y�c�׳�	�d�1���b�����Z�/I�����&/c���Wa��
 \��;?��	̈́�<�~2��K�5�����o�B�T
䚙��� M��\�qFV��X6��q�~7~u_!��R�曁d���a������~��"c�ܡ�W�4�̧1���d�7�\x;�	�e��q�&��<���/����:xj��͆�~Y"3u�hC�f�1�GҿO���Ņ���SY�����Yy�[��ӂb'�*�Ӊ9M�[~Ht���c���*M$eld��_��'�f ���z�(��]Î2������}���e"��~$��`���O,�ޫs�)e`�}�q<7��B�jX��\\7�vz� �I�'��T�߈��7�.&3@d"���!S��-���]�*�c$c}y�`��@ǐg�A&�Zn/3��I-�z���M�8�[�+3�������4����Iyk���|��+��.ԁ�aL�L����m�{&�˝:@�`	)o:�P�Ho�o|L��
��J]��dU���͹�_f����u���}VD��(�Y�-ϼ�h;I'ȥ�Nr�K���i���_�*��[C��$�=���|뿆n��F�G茜V���?� 1~���;%U�y�����L�o�7����8A��J���0"�M��⮘�1^T�UB�HY�c��X��gX���οe�e�L�5��v{�Ty���|��:?�"5yy��0y�����Ô�I�����I�,�^q�nQ�MHQ��N�K"�_�U9����d�0��,��		`�46m5f�����n'NT�C�k�����Q_�.���nKp·*�_U5|t�W��RM~���!U�aQ,��w��I�3a�wC��z�b7q�i�VK�{ۇ	��2�%�2B𛨙ͧ�-u3*�L���C��l����Sc�~XAt��o��2 ��W�x+�����M����,0"�k��s��ニ�ݔ�ʺO�����$�vHKn��x#�c�L���|D�S�Žp�[|�V�D�Ka��_�0;�)�;�_PKS�q�!  �"  PK  ў,J               11.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��U�6kh,�b�����켨sZ.����K!u��e�^����w:6�����{7'Ok{l�MY��o�����|S����ﺪ�v����Hxġ.�Lx0��ß~V=�vb�����N���~��)�nf�by�w�r��������3l���/'s:������J����q`	ċ���O9^�L��$����;�k�?^��u�7�1+��6u����gط�?CPV�t����]�~���a<gQ�v �Ƣ|�<Of٦��j���h�K�{��Z�w��i�t�'^�t���ŏ�?����4h�I[&�ui�u %�Mi�m=�'��"���i�uK�r�\�6�B����&���Lό���y��z���;������x�c�#�&^�V����Z+z���ӝ�M�2i�&����|fR��)	k<v�+�d��P��_ً�@W�BI>1}O�@����M��ӥ�3�>v�Ӻ���kt\��L����̢U��7B']=���1��܋g��[����u�4���}��viM�N�����G���C��-t|g���_���*r�꽛����u�g.�����FY;����V�\�4�a�W�~k�V{�/ї6M�u����υo����6Ѳݿ�����������7s]��{���N��p�������RQvޛ'/���V�p'I6���i���>�$LpLI�����:�s��$^<�Ei×�ӷ��8'gƷ�Bǿ�}J������^�4�z����K֞y��h���7PK�g���  �  PK  ў,J               11.vec�U�A�������Cp���������y �(�����pS��Hy�<������)AɔE)�4e(K9�S��T���Y��T�:5�I-j�u̺ԣ>hH#�$�GS��iAKZњ6����ٞt���BW�e)����{ҋ���/�(�Q��o�<��a(��F�7Jo�<���c<��$&gy1�w��Ә�f2���an�����X�"���,cy��z+�U�fkY�z6�Qo��fy[��vv��]��ۓ"�����r���hq,�q�'9�i�p�s�ϊ��E����U�q����ƭ�����r��<�!�x윟�=������y�[�w�{>�O|�_�f�ww�#���/~�'+�PK�{ݘo  �  PK  ў,J               12.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��U�6kh,�b�����x�_x{�(�����]��Txb#��3��-�)����q��/��U�����;�۠�ﴝ��Q�,�4�:&�ʀ�������/rm����]g��8Y?��-��[��}�t����.���/�||��6{O��s���يM]K]E�a��v�L����3�x�߬�}~�e7<���"�Yl[� ������L�{��_��.����H�t]�*�K��o矿S��?C?���{�~������?Û���gi�L����ϿFn��G��9�\��ٞ̆+u]a��X�s	L����W�>�kc��G[{��L��U4��C��GU>
��?�q��њ��'�Ϗk�k�������xo��1���W�&a��˳�{o�-��na3�oީk<��L�ۈNJ;$m�����|�-!��4	e*�m����Cۿ���<��\ȭ �R�)n�/�������9�/�rcV�V�%��lw�NyWj�?���c]b�'��?��ϰ6"��c����c�V��_f�0|�M�I�K{ҟj��c+�Z�dP��S���Nد��Rw��΅+kڷL�-�ݰ��E,\ׯ��/zŸ8T�������Ɵ�����Li�����7O�Β�g��c�7�d��U9�k������?����7O��4����^�e�s�Np�}!7�^���=��?(�:��o��)ky��}���ni��F�J169�9W�|x|}�a��Iۍ_,�j�� PK���Ԩ  �  PK  ў,J               12.vec�ՎQ��{�@p6@p�]wwww���upw'��@��,�Y���S}NwD���'C��(I)JS&I��Y��T�"��L�&��fV�5ɣ��C]�g֧iDc�ДfI6��-hI+Zӆ����=̎t�3]�J7��#M��3��{Ӈ���?�g��$��`yC�pF0�Q��o��Xy��D&1�)LM31����3��,f3���c~��z�E,f	KY�rV�2��*���ֲ��l`#�ج�Eo�����`'�(`7{��&���� �8��r,�8�wB>�)Ns����<�⸘��\�e�p�k\�7�?qK�|����>x�#��O����x�^�׼��;�=��'>�|���#���/~S��PK�o��q  �  PK  ў,J               13.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��U�6kh,�b����sy?{Q�|~�y�z��������������a�u߇��,�J����:��������/�U;��a�
��=i��l��/u��ta������ɫG�[�%���#�3�Ա�;�?C�ue�oU�i\L�����x�̜�I�o�6��c+	t�ct	��ٮu���QE���r?����/3�|��v�_��[\׹�3.�<~eſ���߿����M�G|$�^t]�*�K�i\�9�~ZŇ���k+�$�K��R_���[ԁ�2���\}�_Iy�u�w�����k��u��L�Ƣ-��4�a�ݧ�N�Ptq������ڽrx���D��n����'�N��2IYdZ���ePǟ�IkY����x�|�f�ΌE]	"���x�bk9U����;TCŋ72hH�\��5��cé���Q�G��g%ni�.:��Գ�wGQUٟ��:O��X��˙KcQ������O�M�/�ZvU/��g�2���w��KuXz�����_�k�G5�z� v|k���ݩ����W+�0VH�����njw�d,۫���O�l���_Z��h�v�6��,����hI�x�}���Pq��[�:���l��{��6�����b��v�1�U�u�J�������N=�����9�����n���y��!k>���׫�ϰ/{�}�mR��)�n�=?���SQvޛg�e�i�����ϗ:��?�!��_\]m�u�ц�O�d�ߵ���e�S�������n�Ӟ��
g
=o̵�T�_fϤu�g����"!"��o PK�����     PK  ў,J               13.vec�U�a�� �Bp�@p���������y �(2i��}��J��H���e�R@������2fY�Q�
R�JTN2QŬJ5�S��Ԣ6uܪk֣>(�!�hL�$M�f4�-iEk��֞vf{:БNt�]�&�]��ܓ^��}�G1��IH�(b0C�0�3�����-�a,��&2��i&��;U��tf0�Y�fs�l�ӛ//`!�X�����i.V譔W��5�e���F�Mz��-le���Nv�[o���+�c?8�!s��iı$�����9�Y�q>����(_�2W��5�s��z��-��.����������3�󂗼�5ox��;�=��'>�|K��ݛ��4~���I�� PKl�&p  �  PK  ў,J               14.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��U�6kh,�b����s�������&��?���7WO��9-���?æ������������	k�;N�|������[O�F����X��U$Ё���\�Qzb��2����3|}��ݤ�7[�ۗ�����1{��4k�nN;}�h�5κ�̖@�lgXԥ�3g{�oze��y�z.�o������o�n����`����۟��?���V��b=�t��/�-wi,�J���g%�gڵw���6M>��������R�H�O�>�D�5h�L��kO�)m,�+�x���*��*�3f.0����Iw�ۙ&��lZ�����~�A״ϡ��v{�~jt��$éy�m����ف��e�.m[��+A$Еa�\���� x��taf��In�>��))���|6/B��Ma��[�N��'���w-�.T���V����{:)JcђDW� F1�ǜ����e����y�؁�����6�(�H������,ՐA��r�sfm_�ݬ&P��ӖIn�GD�<x���~jʑ6���2��X�����+M���]`.?7:#��!�~����?|�=2?C����s�S��}����g��>��8�|�6?��~E4EE������_�y�0%�$u����e��j��gP�����a������1��?u]������Xj���<NO�&��tzG�|��m��=���uZ��C���Y���X���຾�ƿk�TwU�9��,>]���컪�ESE�� PKI$ٸ�  �  PK  ў,J               14.vec��n�3��@p�!8w(ww���R�ݡ��wE�a����;s���$��O�r�R�Ҕ�l��dy*P�JT�
U��d���AMjQ�:ԥ��j ҈�4�)�hN�Z�V��miG{:��{:��t�+��Nz�+M��]�/��OH>�J���1D�0�3���b4c�o��8}<��$&3��LK31���Lf1�9�e�Y���B�E�b�P�R����L���n�����c=��&6�m�۪oc;;��.
��w�&���� �8��r,�8�d�~�S��g9�y.���%�2W�J׸�n�ݲ����.����Ǿ����3�󂗼�5oxk�N����g��oiq|��~D?�8~���IK�PK�{Q�r  �  PK  ў,J               15.i��eTPר�n	A��AB$�Cb ��K:�;���nf��F:�F�A`>�o��s�{����:�<g�u�y� $Jr�r 4t  �i�����8�X�888xx����D��Tdω�i�At��@ ==#�F��������"".�+������M����	)��(y__��?�c�M���� @'E� E{���Ή��������������O�T�@@G��@������|�>���Xd�x���k��0������2J�tSh�:e�p��񒒊��5�V6~A!a�w�ed�����ut��-��ml��<<��}|��C�����������=-=������������������gOo_���������������������߽���˫��w��B`����?r�>q�cbb`�����?��X�x�ɤ4p�ݞ3��K���t�1�i�RX����Ŀ�|���&����"�_`��k	@����<R pV���n�I�)W�3�ۇ�L#��*�9J��I�Tk:Q��镻�d�b�lA!����6��C���bZ1r�h���z{Z��f�3�$_ �1��և�'ĊΏ ��<3܌8� ڇ�1z��=�A��qd��<�����zV�*�4�O�R� �p�ۏ%Ϡ�K��1S�E���y�@ v]
�w�H��H�"�՚�]8&4�n��Kv��@9l�}�k^� �%���^`6:�o��Gd+(7��_+��4G��P�__��I㒡NP%ퟑ�o�r��Ka���+�~���x����2�D��5�e��J�t�̷J�ab�����l2�J��y�)c����w�s���i�RCSt���R]r�.,�sz�3F���ֈ�=>X�Ҽ<;�I��Q]P�5�GlZ���wmH�;į��O�;�Y����M2�������Cf�zB=�Ӷ�@�ٲ7��2Q#�*��`c�+d��qS�s��"��x�
�cg��S��H"u���t�O�*�+��t�#�-�H��a|�X��#SS�k⁭63Ak��*u\8���e<fs�[YSv~+�`�JJ��B1`?[N����l]�+G�)A�gȊ����@�_���Q���� �$���\�o�����z��&2���
.�����^�7��<�g@ð�4�ó\ZE�몭��Η{c֕$��������3�vf�i�u�7ë `��U�蹪�(�ߌ�}�������y|�RY�N�`�-l`<9����`z,:?S��`��(!z�/��7�3�:��d�!S�Z�6L���x���[�u��W���<�"�Ձ!�ǑA-�jR�8'�h��8'S��LkL �^,����-�?ۯ86$�p�'��&)n�7X�]��j1�֪-���;}�;�z�t�_?1�\Ѓ��aw<__�3�K*`簪���S��w�^��Hx�|9b�(�Jo\��pEz;ϓ�ϻ��݃u�9�@��~i��#:���X�z�C�.��R���cV��؜�G�mj4�q9"�]jK�@mr
{�"m�W��ݸ�Pv'�����pA�U�gCjG�� �s۬.��:���������=�p-v �p*�\+:&��}�����i��P�A��OБQ�I���B���K��&ؿ��ᅯ���'�#:}(��&q�EI�Ų��M�F�A���L�P�uVbԓ!h7�6����}�Ǒ�rj�:�I����M7�D��c����k[�;��f�/��Kl�]�ͲXz��7��I�E�+E&A�q=��wt}F2M�!���8%������>� ��VXr�o�?����*W��G�b^����-�_�[�M1y@˔��7[E�UC�p=P���53]}�Z��B�B�ӗ��>!����&kx���&��ӛ؍x1�W�k�1�2\V����nc|`_�};A��/z8���嬱�7����ZU\r �Q���_��Ї�j��9��	,���]�G-��#���@X�T�I��j{�)���E��"|��p�9j��Y��Q���kr���ٖ@�+���J�ݕ�HzU��,P�]�|�A�IU�SK���r��uft��^D����AX(�8<M�~�ÎaE*�4-��v��Xc���c۴�1��Su��'�=��eW˓�s-1��Q2��.$'�r��~k[�W��$�tX����M,���/��oet��^�mK�e66԰j��8���y��
^���;90��q#:]Y6�]+Ɩ�
d���>֫��ʓd{��tf�L!�o�j���?ң�kY�k��!u�n�;�g�(?�&��)sk���ޕy�e<V��c���R���<%)��f��e�P�>>���`�Q����Z�x�G k��b�{�Gza����{�����h�� ��=N�4��΂�8�FG��]��3z�0>�T8�M{S��P��w5��*�T3��p�t��հ�Q�I�Ũ��lXJ�<M"{5
흍�1[���@�`���^����`WV�\qZQ�9[؟j�O��o�g=��5B�G�;%{:N�L:q�(�5+�X��e �R����L���J�y9�w���2�V��,�'۪�J��ѤE��V��m߆'c���`<��9�[�2-
��<�|@��IZqv	���N��ea�{�Oť<�9I�����[��,�XNap8�K�G��C_;�U�1����>�Xh�����ºn<nO.~h�<P�'����"��aKKOZnv�=��4j�|�e���+`*�!���Nh�*?:�Ȗ�n?r�5��׏��\���P� `d�\ns�5�@��}��6��ߏ,y-i��a�mn�(cQ����q ���X;��P~S�?5�ZQ_��X��U��)¥w�~�L5�~���8��p�%���D7߃9��я�J�8���2��"E���_�^;�a39�4����a�}/��Y}��H�|��".���P,'�f�<��{`�zɋqӖn� ��:�g[�==w ���5����6�=��������V�W>��#������G�{3��N��9���,�����2�P���j\v��A���p[>�E@\�7ܰ
��7�K����@6�|�Æ������?{��i���Q?+2��A~0 j/��P�1>&/*oQ���������n΁I���# [a_�a��k( �{�0n�}a���x ?X��H���[��3���F� 8�$Q�R�>�������Q,���,�s��*MI���y�G���v;�N�_
������m��ݘ�F캉s����^ܭNQ�%_�Q�D��h0f�#�*��Ѡi����7��F�"����>D3:3uC�����[�%��|ׅ�{wZ+q���+����C<c�H��6�Ն&�y���/4M�@�-7{�<�D�L����
���A�e�e�P�k���~HCGl�aF�����i�,ލc�2avf� �D~[P��K���i�w�T�[��B~]��ť}�a����3���<�=��٧h�(;�L�@�5�hP�Df�w�Ƕ(C��ı���G�^�y�ޢ�=&?�5���x@�<O<�p`�ۨ=�<��"�!�F��Z���}�]*�+*��މjq�-bJ88)�g��̙�M��%Lo�cS+��QXQ�L���r\�+�*,�!�qK��u���/ 8�%� 8�@|����V���w��UKHl��Ա����%6��\�h
�-N�2Q�4:iu՞;�m�Ebf����q���l\{��;�F��+�3�M>,�غX��З-%JAC�$� ��R3T� s���QTT܂e�Q�$r�Ӱ���l��:��?�Ζ]�lF=�@ZF��s��Cv�P?3��E��gg'�B��{�ɳ�+�/��;�����v��L�o�����:�8����)Q�x���/�V*gs�������9e9{�؟oY���#�
g֒Nۉ�#^
��R�D��.F�J�Y��M�����b�~��~��j�g�S8����6W�ֶ$�%G
]ۼ��tN��/������8�:�+��b���D{VYl}�nk�'��фeB\2-`���UR��π� S	8­yU�Ф������J8.G��]Ҳ6XX4��H�?����.jO=�/��H���S�+ݚ�p��_P���;y�����O��`&���I$���y,4��x�^<[��Z�@f<>m��Y��
�KԴѡ=_ۤw�'ҤZ��%���Ḋ�p{�T����e�`�0Z�o��%�i=��zZ��E^�Ko�<>z�~�K�O	�q�O����Op̱k���}�Lm���~8U���'�J<J �ϣ^"m�Ng�l����Wx+`V�y���-F��x���!=��WG�q%`Pse@,דi���!-,p�O9��l�컩C�X�/�#���U)^�F���[r�Ңi�fS�|;e��<�G1�� _�g�ҹ(x�j�~���dl޺E|&0�B���i��$���֤!�g����/A�z̥5�]LdL�`��Ӵ�~1�7��d�}�����qq��[�~�:,Vvcf[�L�:m�Q�%�+s|Q���G�$?2���|V�0�.$�������m �sC+Nπ�`�4�E��1/(��l)��n��3æ<�c��W�;�$5��m��q~F��_�����;؆�p8�����@�������Ũ"KKa��
fh��nbD%�u�g���9S5첔=Erޡ;�9��w�������9ɻ��t��@s�!ǜ}C���U�rψ��K��{I꯫h�!-͵���f71�Eïfr��۪��FF�)�J�g��bs�W�'5�v⮐���_��/��t�� |���U�*�C*�hth��\	g�����Q��Md-]�[,;��xΞ��ʚD/��%XQ�{��7�� ��F�7/ӺѲ�[կ�0XDz�]��<�x��,�h-���8+�.gb}PDDA�4x��|'�c�<㩎ɽM�ͨ������6�󗘠_5�S�]���U?��?|�w������QT�*�<�G�����Ȏ��RAs���
@�ǅ��T<�l���/?g��tn��c?�!ߧ'j9��4�F���ӱk������E�?P�%�JH{?�g��^�.a�i�O|ri��"��#���h�~�w��_t�=�*�O��$r�X�ੋ.�肼�D;���q5�Fx�]�����:��o��2>��K2��Z��۸!�A}������_�dB�X+B(�B$�M��>Z�����e�o�$�,p5�&�Β݃pPl����KYXi��d�"巵*���үkak��G.��Ū:��e_����o>�6�9�(�f��d�=떳i����X9wWIT�sݕ����U�a�����m(�v�v��U?�b�my{vÒo�̻�m�/��0��S�I�'��	��wV�:�_�<|�ט	��H9C|����K޾�������MC�U^9��^�y@b�~��y�B�4gɣ{�k�a�������̊�g����!��+h�<��2�+� ����C�F����W�>o�ǭ6��+(h�E�{y�͞�;�a���,y�'F��ﶝne[����m�f.*9�C�IN���n?�c����
��s����
7D3�~�\��5�ۘʵ�B
�&,,V��n4e6	+�讚
��t��'V�\���=y L#�
Gt�9�l6
�'Q%�o�o+��e���0Q�(���<�E��Y�q�V�]&�X��m�H��.��ɭs����
����ǖ�j'|���AK��}!�u�E�kr
��L(��W;mj�*���ƭ��oA<�p��^d�>���aG��̍���YFO`�!R��jq��*^md:�%�eO�k��JC�%b����iMN���f���M۰��%��O=�@m=2�!1x�"eH�a,���R�㗝4K��q���^����1��0�'6�k����
#���P�K9k��i�O՘��<S��`8G�!v1�3 D(�%���b�OCf���y���gP�]Q�oa~�Mx4�u&��Db?\�?��i�����I����u�cm�.���Ǫ}�!���b���ԏ�oH����@�
���Rv>y\���8!�8�~o�!�HV�<�-�%�6�3��!C^�5�7��f��G������ӌ�H����)�<�h�7C����S�V�_���y��J�{\��#'�zr��,E���݌3�n<J3|�}��1� �q��ΰ&&��M5�K |13�)��
/t�?	6�P{c9�9"�3B1Y9).R$�}��"^���k��~`���0�sM�鞧2��-j�e9c��SA��\Ś��,g�Y���=#�D7�������0�DC����0�o��o`>�@�Rf���y��<���hA�u7y!�����v.���5���F�xr��?�NΞ^]�&FK�ߊ?�4��
@�C_3�ڠ���u޽��o�V�*t�j8W�*�vZ��]rA~j0k=
�JFl�7�Etc�2L���$v�܈����E?��Ix�����1/����+�MS��b�ɋC	�G>�*o`�q���h �]F~G<M�퉲1�<r��]����Ag�[A��L�Ƶ�_)W�9�=Ӭ�N7ꭨ��{����.��#�;a+�jm�4r�9�g�K�pR��s�k�w�8O����3��_�;�9���iv���J��U9+�9r�@h�KY��]�%_��Z� ��l���[꿎�L�]�/ӆʷr��uƕ,X���7���g)�~�m����o��,G�����x���G��C	C�����=�wz��O��P9VAx�5��
�̘��nr��$U�PM���⏤�B�<W�.+�?[���R�������-o�l�N_��=�������u��j=�b5��6��"�s^V��Gk�%C�	{��9�<��d%��Y����	W)j�S�5א�%H'�f�sYT��m��'(#-)���W�7:���|u�v��o���[���$���BxD����"��]ow�)�����B�V���{�[��Ul�C)6�I jn���xgӮ���	E?zh9�f��ɟ�>�������u	�9�1R������/u5�9֮��yJ�(�p�jh'r13�K�td�箬���!��
���'D�X-Ȯ�#�G�O>ѓ�}��[,�_i���N�J[wD=�b{O�]���Ѳv	�᱂n��Y)�N�&�jɻ�4k�^�4�'�Pp=1���G����(q90�j,�%[&ċV�� �3��?s�|8�Nҿ��*Gq����4��3zܧ�Rf��?�}�e��/cS�nW���t�J������B�5�h�ٸ+�y�JwNv�B�c����i�����TK��n��G�"��Cè�]��^t�>��7PA��� �W.VS��08g���d�Wr~�����.؈0���7�/�p[�wpm@_�\�?w^�R��梕-/p~�pc��><vC!��0p�*�xH~WA-�)@^ɽ0��%��u��D����{F�9)��
�5�r@�[X}M2��`f߉�|�����\�r<��W�E��ޖF"l5��, /xT��m�DgG�'G	 }ٗ��31-�f�X*
(+RgN^y��=Sg�&�ǅd�u8��|n2#��Sz��jP/��H$M��u��_��R�q#2 U�k�Aт	
J4�EA��pq@|��G�F����_/��<������,$$���L�j���?��W-�4��C�,� ��Y�|v.���1��~3��x�ؘ��w����CJ��/�m]�{	ح]�)L��w|C�~Na�"��7�¤���i�U�y�Rg���~��ǉd#�0�_�KEK��T��^z�R����^P�����J�e��FF0?�y�ToF�Dq�2�y�Ջ�(�zƫv�~i�8>1kS�nu�r/T��.��U���m|�V��Ұ����&�h�0�9��.D~W�j�b�[eeG��_m����W�zh�`�~H�v���ѳ��<��/eI0fh����K�vϣ��Z�bI��Q�rqv�SH�����`0�����Xč4Hm� X.)��sC������D�W��mT�9�DG'�|zx�k	�h��Vun�o�
�"̸lq�ntT���E��~PɈ�%���m���>�M�9��r�b���`�NL��{B+.q15-�n��g�[�SSjwG��{�w��L�-me5����\���Jy��
߰N2v��t�$���Ԇq�3�J�띵�]�%HL���ɘ��%F_�r���/�P�I�$XVT�Ȁ\��4�D1���Z��X:����(�������ΊR�ܸ�A�_M�O�wXˆ�Ž�<��<w�y�#8�>�\����=LZ�*�\1nr�>�G���D�=^t���U�{(��xg������]���x�1J�VI��6�|�����w��3�W��y����+���^b�0�a�]� X�zm~�q<±\*6U!T@���Y㾲��� wΔ��є̄����$sv]�DrT�l������=ɮ�R}��+����)�@�������!�:�|�X<��"����/�ҿ��ચ�5�-���(Ysm��"����PK��B�"  �"  PK  ў,J               16.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��Y�6kh,�b����s��=����sA�7��v�w2�o�7����5��������Y�T�cձ�m���o���4kփ�-�����"�0�Ƃ+o�ܭ��~�C�����rsN&���!u�=��{5���8��aÿR���9�@rk���b+	t�at	��ٞ��m�������v�GY���߿���e��o��,��3�k�~��Vm��?ækޏ��ui�u F�kǬc�{[����}Z�f�f_��3���㘩��IÉe[�Z�����}���zWw���LW��B��ve߭�'"B�34l|�3T�����	���=�Z�6��;ˢ�Y�5|Gw=����U�)'V��3tm:�*��:�G4�}fa���9�,�ni��]o�퓊㖟�۞��f��c��=eW�� �+R�����{�V$0(�@�ĚX{��7��|�p��Ma�)�~���EN_	w|�-�{��'1�ܞ�-ϴ��u{�`��{�m<��!Sr�ʿ��6O�{����R]~�K����ǧ�X���/֙*/s�dU��O��b'J	���)�}8�����E��Y���������#>7�	x���n�vu������K�߽=Pg+�����_���\"?�gx.��շ��湋�"��^����8\$�˽�{�L�/k�8��e�y�Z%T����$=�����=1M�'<���<y'���ٌ�����Ū��� PK��R�  �  PK  ў,J               16.vec�U�QЯgv��l���������/�.��;���%�!��������$��O�,y�(AIJQ:�FY�r���De�$��*�Q��S�ZԦ�wՕ��O҈�4��s��洠%�hM���9�e:҉�t�+���7�I=�^��}�G0�n��`}C�pF0�Q�N31&������	Ld����4��o�>���b6s��<�y��n����,a)�X�
V��Xe�Z_�Zֱ�ld���mշ���d��CA��^߱O��r���(�҈�I.N�'9�i�p�s��BZ�.�\�
W��unp���m�w��}�G<v�'vO�g<�/y�k��ַ�����G>�/|図���?"��Q��o���� PK���s  �  PK  ў,J               17.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��Y�6kh,�b����g�4��]�v\��X����E���5:�M����k�ۗ���V��_���!52^�D����)�nfO�zp�R��X�@W|�t��K�͟],]���M�W���FU�e-o_�Y��M"�YI��[���߯9�`2��5����<{���S��|��v�A�FC���_�����q�����う�ȓY��w�XŌ����~\ݶc˷p�T?�<�*��U$�;�p��?I'1���;��6{=��ﴍ��s�'_\���b���e9-S���D�s8�Jc��Ύ�(#��?ô���������9�u�������C��4}��YO�+���l�4wX�H�C'3�U�a�h��nx\}ڛp�wgs�ޛ��>Se}��AA��1mO�_6��nZ�[oN��k����Iזm	 ׾�#�&���8�ʾ�gx��/�ze��?�vs����SO3���<c�{���O��G��{\���s�S�mG��K��m��W������]O��w��;�Ϥ풜���/gp��ί*�?�՞��+�&n���I߂���?��:�sc��'�֙�� !���|қ�/�Ҝpy�Ե�jN�ڂ��M�����3����������}�1��ucR�n�Q�ç�|3sr�?K��ͺ�HqK�k���� PK�� �U  �  PK  ў,J               17.vec�eoa�go{���@p�]�����kqw-��j�r��d���]�H��e�!�,%(I)J'�(#�R��T�"��L���թA5�Em�W]Y��4�!�hL�:��lNZҊִ�-��^v�#��L�ҍ��葤�S�Eo�З~�'�v��}�!r(��F2*���$b�>�q�g��d��91��Mӧ3���b6s�˼47��-����,a)�XΊ4+�V�Y�Zֱ�ld��f�-�V����d�)H#�x���>�s���0G8jw,��q�'9�i�p�s�O���E��)�
W��un�ݴ����w��}�Gi���Oy�s^�W��w}+��|����Wg}�o�G?�(~�_��OZ�PK�@�cr  �  PK  ў,J               18.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��Y�6kh,�b������ѩ���������;s�H���yG��?޺��ϩ]gN��v��D�?��v���"�u���-:��x�.�L]�a����3n�5h<�tq����RW��(����wڪ��2_�M�Qq���5O�e����[79��2�g/u� d���.�c��ܿ2�y���k�߭�;m���Y���=�h�����ҏ�������oQGk
ي���0����,��|<)�~����	U��wʟ�-�n�n��7UEQ�i����°�)F�-O����W2k��&��2��9qN�K%��[2OG>��~n�ʚK:��'�<� i���r��?���gu,�xRe~��c�����su�)�N^���9�䨗koF���V=��� iK���6��^i(9/*���k˺��+�uiqqi,j �eo�T���Ly�q����gh��O6-�l�ߌ�)�4����m�����>s�O��Ɨ��VJ/�w���D���g�5�L�4�T{c��	�9�J�(��MjRe{�B���Z�_�ɛd�g���� B>��~m��=��'��Ĵ<_U\�r��4Q�@ǅ335�r<h������b^�W�l;�s��vN�|ú4�|�Ru��q���6YRsj�:㗟�bں��bƢ���o PK��B  �  PK  ў,J               18.vec�U��3_�؊�؊�؝���������n�[A�Q���6�&"I���!K�<E(J1�'�(!KR�Ҕ�,�(Ow*�JT�
U�FujPӦ��M�R��4�!��L4�MhJ3�ӂ����;md[�ўt����'�����w�=�Eo�P@_�~I��d��P�1<�Ĉ$b�>�ьa,��&�٘��&�S��4�3���bv��9vs�y�gY�b��4��2���
V��լa-�Xo��n����la+���v��|�n}{��~p�C�;���~���$�8�Φ�q.��y���e�p�k\����M����]�q�<L�xd�X�S�����}���w����g���տ�i|���!��i�PK���p  �  PK  ў,J               19.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��Y�6kh,�b�����:���[+�V�_���!U�\�������>�gXpmZc��ۺ�[g]�����s����i��N�g�t]'tu�e�Ƣ]�lzec_�����������|���6{O�oQ��m߷���W����s�3�F~<y�[���f_%����XKЂ{�O�;�WJ����T������[�wڪ��WW6����P� �o��c�����w�g����O���Ƣ���4�a�1�5'�_��˵�����WY�g��m��4�ㆽIJ�}u�KKwO�)��\����c���q�N����:��R�'�Z��e&�M5�åAE^���LQ������<�?�6�H��r0����*�R&��L\�F�(&�Z���A�0K*�z�?Z�+�.Xa�ל�����s��O>ˍ����Y��䰭��ӗ;�_[Po��t��O]i؍3:��.y���X�������"���{+!���A��O�#��4~<�|ej��׾�5жО�� �}�ʕ~4���X�Y��)����d/���єȥwVY/^���f���|=G~i�t�J�����_�<�E�ͭ�ԥ�����M PK��]��  _  PK  ў,J               19.vec�e�UQ��ܙ�b+�b+�bw�����������	���Gk}X��aG$I��2�O�"�œL��%)Ei�P�r���s*�JT�
U�FujP�9�dm�P�zԧid�X6�)�hNZҊ��j#�Ҏ�t�#��L��ItMr�M�Nzҋ�����v��4��� 3��cx�����b4c�8�3��i^L���Oa*Ә�f2��i~̱���c>��B���,ai��ev���d�Y�Zֱ�n��F}���V����L#v%��=�e�9�Aq��H����1�s����4g8�ƹ$?����%.s��\�����oq�;���y��4�Gv��'<��y�K^��{��o�w����g���y�2��i����)�?i�PK�M5�v     PK  ў,J               20.i��g8�]�;z�-�{-z�D�(�ED��;�3�ޢ�3$�N��Q�w�3���y��|9�9k�׾�u��k��B�A���+�)00 ��@/���x�8�xxx��D��DO�ѐS�R2�212���3��s2����s���a└�z�/,"��!DO������X�Y��?�@��!���``�a`�a�{L�����?�������S &&66��7���&�!g�ǥб�cu�
I,�gS����}�.������4�/88�^r����KHJ)�QRVQUS�����-��ml?��{xzy�������GDFE�$%����gdf+)-+�hhl�7��"�~����ONM�����_X[��������?=;�����A��ǅ�������E�ȅ��������ȰqXq��u�,�(X�B�)�	؄uO�>��&|�.����?��I�����/���� DX���" g�)d���q�u56�Dū����Ͽ��Bn�h�����}$*�`IeC�/�P�z�?+��qTw8c zN�z.���8�z��/�*�?_qaz9������w�����됣��ݗ��<���X�����ԕ�hd �a�Cry�;��!�o�6�;x�rRwD�E�{픃�8���a����#�y����#"�kT�Iu�B�U�Gy�O����A4@jM$����T����e7p9g[Ef�R�s�7;~/�2@`*�F���[F����ꔱ�!8p�e��)���:Ŗo�LQ���x\����x��������.o"�;����{p�F��-_s=gf��SvƢ2T
��]��H��Z7��ۤ>�i�}��@e��g��d4���[��Y�*�q��� >%��.��,���?'�9΄n�ܡ�TBP�C���;x�Ájgͨ�������,��5���{h����|���nW��r�}��j���/u	�J��Rr;P��/5�>���-b���R'�;���<����=�{�}�RVG�Oݖ�J�O�˔r��� ���on_�d���M�#C��0g�ډ3M��f���]Ǒ���[�r����!�#n�}'�e��`��lJ�KPw5�v�P ���-�kP)x$��e�4��+F�_r>���h� w� �>��Uv׃������.x�P�H��LG��τۦ����܋mO�
vk�v����k=�؝X6��]N(H;�X^�'kE��W'��ק��J�h�,�@<�m�!��󥠰ԪS��{^�(ߴ/q�[�w�Q⫖���QoFx��]�h}O�yL
#�����r���q"�v*"���/Wc }��T�f����'���1��҅�9�FR0���Q^|����#�������ײ��L/\|р�W���,�L�eY?�yJ��)��;a�wl�~&<��o|�������r!3
��{4xm5&��'�ko�7_� 6�Kja6o�M��R.�D"����V�W!���u��=�q��NJ/�`g������1ò�9��`��5>���М^Qxc�!]�&M}eI\v�zHv�ć���J4<�����>[�\��;�$<��\�bPUL���[��'�����Y�4L�S��y>���;��!��/��t��ѐ8�Ek<��Qo��	��__��d6�o���é���g�MB1�ե@�4�mv�3���k�n�	���p%Q\=L��"��Oݽ]Q��1.e"	���x��0�!���3�0�J치�RG^o�s����وX���n(�8
1�?�/��#<���/�J��1k���*��������n��o�'�����4��5�A�� !�J�| Dy4�&Q�2g�ِ1k�2���֜�a���*��>RA���Y�`���.O�G�D���a�-I�.R	Z�f�o�f�؟��i}M�����*<O��6O~jM�S҇���z'���+�z�O�UQ'(��\OY6�f쫥�1ė��C��T��h©�5$e��q�,�B����G�d7�G���4�͵^9�
B����o�[IX�D �0� ���~٦Aذ�	;ᗁ�k�ɒ#��5%)�0��JFʀ	����Xi��k!~v�!n��Vv��U��i����l\��}��υ\����������T�������3%^ݰ�,GK��'�|k5)�M�(�)F��1�l�Y(�@��%�[�/B	+4o2�u��ȕH�������H��Ԛ.����y#�ԙ7���������HN�d9&AUX/&e'���p6�=����e�s��;e�n ʤ�r2�Η#�bO�����,�N��|(����`�D~%8w6�$$��NC��r˨q���
!{�;�MWbB�L1?��IF�,E��@����JmϞf�3�P�a�_�����`ڊ~y�*I��GЊr�po���Cf��,�X�ħt��6��ٚbjz=C=��y�d�g�x�!JNvW�?����\C_��K�6`:��?J7�������ȅ��M��IY�Su^�������_����S~<k��y+����m�ԛ��&=V��C|Co��Oy��Zm��Cҝ�K~y�vAt����t ����<�h ���ŶP&�>D6��c���#M�3�r�//�eazY�#�}�ce��gRy�9����!�$�zY���|�ɘ`;~:U��'��`䉓�/���}E��f���Y��_6���s\F݄�S8{&�×���n�e"iVuƛ�Ŀ�"b"5�=#9�L^(�a���e�KfuqH�מ�ZrPd} h<�����wyJ�??P�_נ��N=�,p>~v�����\l(�LZe�f�F��R���� E���f��2�޴ޗ�qTN�jG� �%��2�����[�۽%�����~�]���U}L@$}�J��ba�@����\o*���xw]0hJ���,���0��O�T�PԸ��¨L9�FI��K��/{e��~:�܌,}s��{��k_G��Ծ�����V��i`H�K~Y���b��ŷi<�� �{3�w�_d����Q��D�P� �����pg��!���Q���N�_wbU(Mu	��ɥZk^�X��:�z���b��P��%�`流H�i;��5����}%�ݡX~Yo� )B��߉�6���čN�։D�jIgN�P�gbxt�r�mb,T��@�G��l�􄕰���O���!���o�&���-G^�7�����+E��3����7���;Z�c�7B���c���u����<���Q��̬����I�c�y�r������?�?�U��	߅�L��"�%4��wDM^��}cU��LA�n*�Y�d�M��b+-Gt#8�5���Y��*���PezV�Ң�؟H���Ǵ)s)|�_5�	�KP{q��
�2�NM9m�ڰ�-��,��JM�����P�� cx�<2���&Uy����R�J��e�h���WW�:ߧ�������r��e�o&&狨��`��H;�34@%J查a5�ݼ̟�l�魄w��\��j�--�`�%���_��}�"�}�t
��5���S���}D��3lb���	x圵����.+�6�t�d�n�����M_:��uUCQ�T�I�$Z�{�g�4�	&a�A�A��8YK��6�.ܰ��{en�� ��u��������S�
&���w����US�Y5e����YN�}&�y�l�3X�B2�g[1�(Ԑ-�_�0�%�kAP�5��?�u���f�~�Ԙem������|qbN�/2�_R$1��t�YMWI#.�q�+S��fTh`9���G_���A��h@�?/�%��5	���m���έrI˰2&@��(����Ni���vU'�4uQ��8s���e�'q����̋��#A!Kb#<e˄1�r�d�uN����Շ��EMu�Oӑa�?8�LpS�1���M��@,{��/�:�)��ܸa���������C-�|�)Y�Fo�:��x��>�����6ݦ��I�K��]c£�����å�~NSy���d��xx��5�&tp�!�e�X��x�D*j�7��m�j��0�!y:C�������UW�U궸6\�糹iLm9X�����p��5��W�_��xRbԖ�P�>����5�u�7鰔�к\x�&����O�Eg��`�5�t17/(���ND^%��N#Z�J7��տ���Y˔cq �~��=�5P���>D���<֧k(��	�8N�L�HMJ�qVJ��ތ��Qi�����ƽk��]��uU�̇�$���"����:�!�^i�𕭜w���u�$���_�4.[�U�o�ʆ���59�h��T[�M�_��=�ДE;Q�a�Ekǆ�%D���Hƛ���=�����Zbu{DU��y2Ry�|�I&���\Peʠ�>'�t8h�@;�iT��b�5��!ܦ܊��h��A&e����͢�q�ol^r�')5! �>��u4:1��\�+��gKl����X2<x�	HgG'��dXɔI�����td�ݯ��f��!j�[���`��kwZ�� d��ٟY�b�GmH��Mn�N#��V��Q6����p��[Xb4-���ٜ���a�$Kk_����tzֺ�zl�����D	�s�]��7]�P4��X�LU��Xn0���Z��V��1�Kz�[]H��XZ��G	!��(��p�e=دTr.3y�;��� e��U�$�Ƹl����֒G�nx2eu[��tr٧��I5�*����z��1/���<��Q��y�������H�
�(��{~����[`'	�ĖV�6�b@��n��(ټ�x��f�q��C�k'�wy���g�ʛ�f��,U�P��*�mZ�"�y�4��%,�5H�)��fi�3W"H��q��&�F�噙-L~Px�8~����Z��R�i%K#	�g�|EˑBN���ZԆO�р�a��8a3;�  �P�� *��*s��]�T��g>���V�ꏚ�D�h�@�n��qi^3J?�`���DQ��%��E�WFEm�m�H�M� �9�,j �DpnOY&բ32(�5
>j�e9�2G��s.�)5���sג��i�����O��6������_-�sNQ��i���+z�����Q��{/_B�~i�L�!�c8PHec�ܨU��z�t�Lj����#�eSl��o����l�����t�u!����N�r����Xd���O�� !b��,��Y�E��chű����M�ʘSQ<h�� }�o�����5%��y_.^`g��`�6Hӿ-��|�{�6�I�����Z����1��Y����#%Wƛ�d�'��N(3�}�,�aT�_��_m~r�,�#���3�KӍuk(h���zx�IF��u���6�!W�U:a�	'z�N��^X�0Q��DJF�\L�q�%��p�պ�Љ����Ā��y*�� 1"��f�×�j�)"���x���0�%G�o��(�.�J9d���I0��9�X���O��g}-m�F�1����{@ �Ƃ��rΰ�X�X�AWh_� ���P�1�(@E�H��!�4t�n֕��`_Ey%��캥h:#����o�:N���D��i�O�x`¡N��U\��~���n��/��8s�]��T����!"�Wr� ���6��y��w6^�v��R��~��py-���H�����;���7Ɉ d����ݕ���ML�x���hQmu�&$���J��}����o;�E_k�u�����=7��Ӟ%�
�C6�<���$5��/�х�J�J�oi;�O�����*:r��c����s��>�.�nYc���H�_��Vud�?MAw�pAR�Vȸz�j�����ӈk���1����1	O�P���uà�%�`*w sn���P��������Nxpm��B`Dj����XL��-{fԌ�}��=����`�8��=��6n1�X$�: <"�3Ya=�l�d؂:���}�J��wOk&y�����&QZ��H��ޯ�e-�������6�}��<:Y�bk^l\4d@�kM�Ӓ�1��l�
���Q���yJu��Jg�pi��P)H;��P"�GL�T�1�H%k�����uU�Q��Iu�x��m�u��OZm������*U�c3)�Y)tp̴�2��e�n����Ǭ����ǮV�a�<���c<5'"IJF�Y�����hxV
5�\Mz��[�?��&/�c��x���׈T�&����(�z�[.������0�:� �E8ʃL.e��E�U��e�DE��i��f��u����~JV�	��B?�w��$^bZ��CWX�?��Xk/�:7N����\�R��-�4�4� ���nz<�Cp�Q�fM��7���&3�{2�x�oH�S�@�?���'u��ޙ�L�[��̽���#�*,���+���d׏�9��]
A�fW�+��������-Ѐ�4`�x�M�NO�GJ\I�l�R�=���AO��
�7z{�]�wɁ7�-���M�J��&��w_z.�g�Y�#���y��Z@��!E�[�X��S��u�0�\�%�$�1_���UL�O��Ջ��a��V�d�n�O[�r��ܽQ��6��+�Ky�<~�&�M^P�iP�F)"�* ��������@���Z������m�6�	����,Q�5��da�s#X�ii�T[�k��(�/����S��+O�%��y�tOO���lau��*m5`A�4���K�ET���h޽���:)c�I���k���_�eM!�]�l1���,���R��	H� ��X�w�Ҕ�����|�ӟ.��LM�)00Gڄ^R��5��VC]o$�A�+!�l\�Ǣr����UY�)4v[d!�ϥg���w���NGͥ^F�KU�����ڂ��'�&��*6�лI�z�����;���A-�K����A��
k�i�R��7�6zwb�
��F��(4��3A��N;����I<�"�����E�?#V����6�7?���y�H>�aD9�/wޮҗ�ٵ�_5O�qC�ۣ�WC�Et)�o���c{��x����P�Y��]��Ru����P���И*@��t��O�%0X�)�6���_i�g��ů2��s�H��nP�����KM�V��09���?�>؄Z'9X�6�Z�C��"�XnWHnhy�Z�]M>Z��Q����H	=�I5Qb��ߍ�?�+��4���h�"��w�����:��(��&��,ʨ�Qc���G�j�ʆA�p�I�r�����e�>.�瑮�lO��j�Y(seXܟ�ibQ�ґ���+@��6����q@�T�B̿J��1�b�rA�U^�:���Q�e��O�� LqHlk?�iہ#N鬗�%(���>W�a�q�E��T���[������z&+�(��ӥ�Q&��_��J��M;�ߣ����)�_�� �J���"!��[ǧ�S��t�+�j��V=^fI@E���j�G���;��V^Ľ_�ė�H�w;Q�1;�]���:���*���,�H0�52�?��N��P���"8)�xh �G mKm�[I�0׈�]�'��Z[a@���q5�_=���e6Ә9 k�8�&����g@��$�5�1h��K_ g�$�7;`nL��? ��;�8R��޾����V��K�������7jF��.?�㇝��N���2�q���W��M>0h�3N�b��������Nt����ޞUDXԑ��2|©/�8?qL��
N�;��K��.W;I�J{�l���	��0LA*i�L�^/cTTx��T?�V�2��ؚ�,F�]�0�Z"��UfEÂ��T��C�7�^�꺇���vε��q�՘�)���A)P|'0tZC@Ƨ���׸�oM|���V���0�I7~� +ﮧB����L�:��Qd��V��Q<����ikD�*�Ѐ<��À�w}"~4#+rL������$u��2w�~_���޷P/�Y��C�K�ev`p�*#Mp�iM :��h�%�S,�=��r�`CJc��[5t�1��d�)�W�����!� 9�F1��\s)�P�#�)��j��kN�\毑rqyC�*��x�:4���Ԍq.ɉ�ft.��~�BԮ��k��� `t_Ժ�� ��w���Vig3)�K];g�|���i./�����x��Bo��Yv�F�����gY����T������տ�K}�Q{32�X�� U�e��$m��Z�py��G]��R�F����ZL��J�D��gCsf�s	1��	�E]��ʿ9��X�$o���\���rxS���g��4p� e�@��C�W2A�a�R�n])h ��(&�ie��N�w��
��;��&k����<\B|�p��9������2�rS�M:/����v�O�����$0�al�d�S+I�K�?��ڞ;�n��9�Oc�v_����\~��$��+�@�J7�>-񈭮̋��%��ܽ�(L_�%�M%iG�zO��f�dgR	�J�����ϋj>���O�H�>Q�f~���zڪ�DQ���r<�Ĳ�� (+o�|�U�L����Y��J�ϤI�\���Ĝ
�m��*��${�7b� j� �+�
���|A,��n�C�ԙ�w{c���d�y=�1 �`�){2d�;�&6�ڱ��U��i����PK|6M"  �"  PK  ў,J               21.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��Y�6kh,�b������]IV�K;��a��?G���mH��f���Y���ߺ��P~���?��5���Nݤ�7[ϊf]g+��Z��*3^�(ʽ>�{ڃ�>U��f���6�Y�i�-j��[�*�/���ʖ�?÷U����7�/-�ϰ�Z���閮"aD]����_O�x],,���)j���7�]��N��|Wd>��S���\�/�������R�L�����.� .�E�0w�������&λ�7�PwG��Uy�oUw��*�S��y��N�dzd�bU�?�����Vi,Z�ԥ� �|���;���*��>_0�:-^���Q����j��_���K�$\���R�U$�a�br�ċ�1BF�����s��LZ�q��ig��ֵQ���=�4�?c�U��g��ސ�&���K)����оj>��ց�|��y��*g�&^���W�����v�c��e�m����Ϳ����)ʻv��[�#x��i����gs�h���������� ��Ɣ盚翌��1�s�������rs�-	;7�̿�����~���i��w	Ȁe���7PK��ɕ�  I  PK  ў,J               21.vec�U�A�o���Cp�!������������> ?je8drR�P��tD���/C�d)BQ�Q<�D	Y�R��e)Gy*8���De�P�jT�5���%kS��ԣ>hH#w5�MhJ3�ӂ������ȶ��=�H':ӥ ��IAtӻ���'��M��Ϯ�� } ���2��H31ҽ��ьa,��&2)͉�vS��Lc:3��,f3'͍�v���,`!�X���,��r��JV��5�e��`�1��&}3[��6�����J#v'��G��>�s���0G�:�~����9�YΥyq��~�K\�
W��un�ݴ����w��}�G�����)�x�^�׼�{�]�����G>�/|�[���La����y�+��͟4?���� PK1�y     PK  ў,J               22.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��.�E�54u1��_���\|u���T����3t��a���{S���v��Rs�����������K�+���t�����1���0���K{	S��|����d��/}�>�;�4�?���E��	_��懝���q��~�]�c���,�3ħ�{��������H���*��U$��eY�9��qc����!��Χي�g�ufқ���=uo����|���)�����M�<�OH6���-	te���8n*�<����5�燈�ߛ,��47G�x���1Pk�n9��!ٍ�S�30�T	��۹r�݃]E�=��7v�v/'��^+i����Fm��O��3G{�n�W���Gs�Ź��q|{ i��%�]EeZJ�	7�����D7D�>�j����y��_�y����:s�s��u֬����j��Uy'<\y�S���L��]�C��u��9�eJ�~}���T��m�	��2�~?[W�:7OW��)����?S��6;Z�c�s��Y�Ɨ_���)z��fo�/Y?��~�\~i��k�j]s�4h'��<�|h��$�{�
�<~'o��"�JcQ�â. f� PK!�Q�  P  PK  ў,J               22.vec�eo��;��!8ww(���������]? ?jK�C6'����N���$/�9����"�œL�pKR�Ҕ�,�(O�$��n%*S��T�:5���D-�6u�K=�Ӏ�4�;��&4��iAKZ�:M��][ݎ�t�#��L��M�[R�uzҋ��!����럤1@d��P�1�i&Fz�(=�1�e��D&�91�n���4�3���b6sҼ�k7O�gY�b���ev��V蕬b5kX�:ֳ�nc�Iof[��vv��]i��$7���c?8�!s$M��1}����9�YΥ�8�=��/r��\�*׸���v��m�p�{��yd��}�S������o�'o�;��|�3_�j�-Sߣ ~D6~F���ğ4�PK9��|z     PK  ў,J               23.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��.�E�54u1��_��=���]/�y�����ik�w��̪�߭��������S�e����H��й���X�����i;/��zp�V��X�@W�8��,w{U��6�X�<�k�/��������Y{7�0��`���?C���jk*��:��:P.[����9WE�]E�`���"�&���h��a_���0���7��3l��~��bu�Æ�����X���漝� �U֪�Zԥ������N�3��b���,��i.:�n�+��z�.~�?�93�C�Z�c#�ߧ�����gй��O_��*�E]�x�b�E��T�W*n�>�2���>K��I;���,�75�}���R�5^��w��J����E0=7ʷ���<!Od�^�QL��m�%�dP%v�C~i1���&7]��*9��D��;�x�J,���,�싐�]���{��0i^��?�r}���5���>�Mq����KX��Wk~}��$�~���.˵6.Բo�n>k�V%Ւ�5{w��	S)S����gu��i��hHL�r�Ҵ)�0�_" �ҁ�T"�ߩ�%��;���T����?�p`p�E�[�H�c��H #���	 PK�g-
�  Z  PK  ў,J               23.vec�e�Q���!8wwX��������-��~ ~�,4�tN�sS���I^$�Y
��Ma�P�bI&��%(I)JS����|�D�"��L�R���H�QӬEm�P�zԧ�id6�	MiFsZВVi����miG{:БNt�˟$�&it��Ӄ���7����}����� 3��cx���;R�h�0�q�g�lLқ,Oa*Ә�f2��i^�ћ+�c>X�"���z����+X�*V����c�ކ$b����la+���v����ny{��~p�CN����Q��9�INq�3�MsqN�|��\�2W��5�;�z7�[��w��}�P���'<��y�K^��ڙ�����|�#�������[���ŏH�'�҂����PK�#_ y     PK  ў,J               24.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��.�E�54u1�����k��l�:�7gS�K����y�O��i�-�ƾ@:�2�׌(3���nf�˙�n����a�u��};��/��^�ԥ����?�1.��c6�{fv��mM>�nٟ2�c��J}"�V'�}��OV�����]�~���a<hA �Ƣ|�|]tڦ��w���g����rO��u��w��N�(���d˿���_�G]���s��]O��3��Y���&+��*3j9	�Sn��)z�%τ[����Au-��;�4�MV<i�a�ok���+N�y�A�f�/�E3XEF���,�K6�U�m5	[�\�u�{k[nߒU����f/۞�͖�+��B[縢G��e�Q5�]���X��*@+�fZZǿ=tR�N�l��o���?Ӟ�\�P���ҔȌ���ʉޟ{�+����{�Y��*E�Zv߰��kTd[iiM����/O��w�M`��N�n����I,�B���q�+M�/��2hWL�1���0��ʵΉ��z�>3-���]��:z��b��.l���sD^�ɚ��V�*K�{��OkkI�]^˴�E�קu�o��
tw,?��	 PK����  I  PK  ў,J               24.vec�e�Q�=�zUl�Vl�����������V�������˸dX�g�as8'")�/C��9
S��K2Q�,AIJQ�2���$*��De�P�jT�F���f-jS��ԣ>hhO#�1MhJ3�ӂ��J�h�Lm䶴�=�H':ӥ ��I�����'��M��Ͼ�z�b0C�0�3"��H�%�fc�x&0�Ii6&�M��2���`&��͜4s����Y�B��%,e��r��JV��5�e�٠�1��$of[��vv��]i��${��c?8�!s$-��z����$�8��r.��y��E.q�+\�׹�o�ݒos����>x�#�������%�xm�w�V~�{>�O|�_��y��Ə��O��ӿ�'��PK��w�v     PK  ў,J               25.i��e\��������V:���;���.AAB@@VJ��VB��n�Ni�������澸��y9g�g�s���f�x�����z `� �@���������Ĕ$�DD�4O�(hA����Ll<`&����/9_��		��bR��<�B�	�E@@@LDLMBB-�L�,��l�N 9>� ����� ��'.���#l\< >!�?��ǀGX�؏p�qqqp�͆�����R0���=ѱ�xQ
D&�g}U�E�;q�&h������3j���`N.!a���b�r�
�J�*�z��F�&��v��o��}|������G�|����%-=�k&,�������������������wOo_��������������������������%������?\X l��i�G.�\�pp�q����z�r\f~<
Y����H|�W��k�XuO�l�'��	�??����߁���"�_`��k@���/y�� (����Q�͍8}�:�"�a����9S(&zU*D#�-��%9s+}�~I1���Rf~�1;��|�KkK��v��BUK�����e ķ�ֿ�`�nE �ӏfK�I�:�	O0�Sr�[���]���s�QM:2]�T.�}��	��h�8�f�Ln}�KP�; �>CӬ�3w�֗:�����~�c~����N/�c ��5����%�4��]Du�'�����7٦��o]U�Ϋ�P���,
�]�I�����c_K�D����l��-p��i	V�0�,
�iME>Txt����e�*�2.�A��=!Z`&�[�P[T� ���Geoeg����]
4�ˡ�~��7�~~�� j'��~^���|�n�� T=��Ql�������E� 1���B��E	筠~154�?�8�ܗW1�]��.��ҍJ���@�=��  ����~Y���Qb�$�8�LKo���t�FነUO�ىEUf�s6�r������Ϡ�]���K�#��u,Ɗ|�c�.
�����dM�ZG��4�Ƹ�ŧ�A��-��EgE�1�4�'��K���opvM�5y&3X�y-�<1��;ti��d<��\���R�pc1�-�<�{����G�Z��aO�^Iԏz� �}b8��>�6�ȹ�S���]��?8:���ڕ����1�g�<l�=i�CB��l����9ֻ�\�,���5�]d�a�F����۷y=���=�A�/�0*x�Q�%����^�A��g��1��M����!v%��`���S����k�F��-]���FE QR\^]��w��ouV#��~2��#����3q��i��?��H����DD=�qhi��R�M�}�o�F�7���8�	�b[qw�Na�=��J�%�`�^����:u��P����n���<��>"B��0.B>��ca�($PO��p��Y���*������̂��s� <���^qI頸}C�^+��j
�W��z�Si?i�m����՞� �/�0�V:�P�.!����������ٲ���z���
y���������U�{C�+�g����w`�E�b�x�>E�����sɽ�r�>\T�8��^��m���2��H���4�#"xWùf`<F[��JH�y���;;��J(�
�h���⾧�є\�_+@�����ۦ�҉��$�(>��/���+Eut�쟷�a��6o9���i�?}e�ʤYA�b7���ڙÞ�U���/Z(�*�v�y��\�«�iR�)^<�F���J����>���mS�u��'d��iR��w� �O�_�1r�4���ڿv�2�)���RsF�U���z!�|:)"8xVt����*��(,���͔{���QS�9��?�����~ M�;�������b�L*<dښ�(w;��G��_��A�,>�3��3Bc#�}=�f�'/zt�yFȴ4]r�Vӄ��c_�r��8�D��p}c1,�!s:^��q���Uޗ�ԘeH�+�;}T�eN[^/�w��h�(�b79��Is�ƶ3�mmk:�<80�0,G^�_�bM�|iXV���� �錚��I�3��������_Y�Zi��V��L���/����*�GoVA3)럏�sY@}SB�JڊSӿ[��U����:;�	M��Q��֏�B�*�~��)g�>ɁDě�O�.��TJT@��o��JT�{S��<[�'���z>q?�CC?��)�ٞ��Fw���l3�P���~��i�B]a@z[���\�`y��B�����r��A��9�c܍��+��6]��0R�F�nfA�qK�8D�i�lp�uٕ#۴l�d�4�\~k�CэA��C���4I�I`�=\X���i�ELX'��
��/�*-�Jb��U��-�|x�\�/nR����5������q������gHf��{M7F��L�<#�A�n���I��.�w��nm�J�;[������2����_%%e�r/��1 �H�č򖃍ȷm��E��}t�Tz��6'�OA�ZZ�d�̒��7>�_*�W!]y���ѝ7�잺��Y��O�U=����x�f[��ͲHP9���ok\��2�s��cX���e�r�|�lSEm1��'�
؏��Ʀ>¾�!���^��"y��qcĆÞ�*EG�%���w��N/��r�..��A��LG�6�c���Cj+4n"Nf<6�H8�co�-�Xe�� �8�}Cf`�T���R(4��k׬� x��T!4��B!A��v`�/k�Ԟ{?=`��Py��G�N�<t�
�j�2e�H��M���U=�16^���tL�˖�k�+	Q6i�J�t�?[mh! }��	����Vlq�\b���7EFSQf����w��Ƿ$,�^�Z�8v�_�x�![~!I�qi��n���Sׅw�}}�]a����3�6�s��^Y����eGzK����:>'���6�tǙx�_��x{�����w?k�Һ���E�S��<p���r1�c$C܄�Ҹ�<��}�5��L�WC��ò��Gvx�9�J�a��'0M�.N6�cb_&5�����7�_�~@6r�M�.���j��rH�l�ю��v�f>��׏�b_B�h��$��{~���L�1F��Wld�B���v4<'ɗ��n��s�ف=:8�3��(��;������C��|?'���dq^__1L��9-�d`5��n���bu��R��l��w��4U:N�78z;�Pz�E_:v��,1[U)Z�dyL�q<Lvm6�B�����giĞP�$��,=�ƽ������w��i=�7�%�h8�F@%k��M�1g�6�~Aw���h<t���Op䶸c�^�oZ��*���4bI��,=c��X�s��1:q����h|������y�Zi<�����G;>d���(ʅ'y��	�ɫ�J��Um������=i�h�#��$W1+7(tOS�G�M����٠fc��Z���Oo�"^} ���}���� �{��F���?:���oߴE�/�:��:��7-�4���,#�Vj䫫Fh݈��f��% ����_�qZ�=��gsȊ���C�թ[����b�h�+}�!U��'7p��Ȫ*���9~5{O�GF�BSm\:j6������W>/�I1���p58��i>##?xN��b���6��G��w �*.���]�����l񠫺a�v��}����	��B�֮����91�yx�ج�����r'6c�NQ�`�|�]h�\e���i�&{#���0*��	��~%��tɢ�����{������vUߢ�'GR�"j�����I.��=th�[�e\C1��w$lѺq�<ĭb�'��ah/%w�Qc�|ˢ�ؼ�p���`8�?��-i���l2���b�������l�r�r�O*썖.:�=CqMy�_��S<9����j<�����&��H�E�4�*�>��Qx?��.�!{�g�"+|\\�C�9�Sg@1�`�'Ӱ<�D�(�����T�΍��f��C�9.����_�n=Ox����{�q���)��&Χ�VF4c��_����Dd�e� ^<y��"�:2��קUF�70M��Uo���nGP���^eO�(S��l�tv֚Cu�������F+����Y����~p���s��'yؤM���&��(T�W�X�y;$ː���Ix$����ϑ[W�B|e�}�W���%|i<�{��e��=ȀJ�eno��)<�\��!M����R-p�-��1��)����fo-�y}Ju��́�VY��s2MIV��u�'.�J��(h����e~��jA����������O��� �M��J%S�h���YCҡ(���X5��"�g)�7�{^��Qu����K0�8'��{<.3H�1>���-]د>1������,,�(-xb�����[_�'@������]���9���'ɓ�7�޸�6[���t�������M�Ei:i,߮�4��q�i��.H��YW@z+�	�A1��lEY</D��}��7O3y?֕�N̓6�j�QF��b����r/�͗%r����O]j�&�����,�l�.Yo�ЌH����m��c�2�7��� ��͒�ޗ�榚�>�	���AS�c���cޝ>
�_�U@��q����AӁ�mj=+|�W��r��;�8PY�\�&�2����l�*%J��ປ4�)�W��2�G�G���� ��I_{������ �B���Ir�Z��"�N� Y)5�Oq�)���\�6�g�|�.�i�Zvo��Z���L���,7�<�h�0�.�o=�V��L��V�����/2ˎ���Ŷ�v�".,��ƵL�򷘯h�W�J�����a93s�9���Bh�;>UI��5��K���?�e�d-�ғn.O '.�Fb;Uv���\�O7g�83	ǒ��<;��2%���z[��B��kْ���c }AP�Cs��̭Nh���U"��o�/N�����M��M�;5+/#��Z�����T��6*΄7{"�����?#ҡ�8�ݳfY	g�����S/��[����U�z��C�,�5��GB�|��[�,��u�4�X{�\�5���Lx].�ӚK$����u��)�"���=o�(�]�w�e]�ZA����~����qr�e�^aI҅��W}�a2�qc��7�e$�+����=������NX���;,� ���L$���Ԡ����\O���/>5�m�~��UͱN6�~��PW������%1��g���
���&�u�i�
�q �;}P�fݕKn�29������,��F��FM����|��
8U�KP�&�.�y�g�7fۂ����m%���)������G�M��S�tI��y� �z��� k���WU���Yۋ?�,/��!�Mw�~"�gh����u�9�e��ܧ�5�wY��x<�K
$�pJx�i.56��>����i�~)��0q_��SYix�<#�������~���e<��)�X��B�Q����l�
����
xp)��*��vۘ�bO�D���<�3�&3��xkq�Y�z����1)2z��ߑ�8����&w���Ϙ}��& �4�Ͽ+-��18N)_�"1���E0�K*�sam@@*�fO�]j\�O� .����eE���O�m!�Y�7Ʀ�s���B5���x���CcA��6�R�42A"�>G���_wF
)O=��Ӥ(�Ї�EL��}�R�/���ŤWg !Q{q۵*�BJm���Y�۩X�*%ʼb���R##o�hߺ߶Za \G�L�s��.Dʑle���5{�g��-zL��cX:\�n��H�aWP��Rǣ��'ì�0��jl�d�ZY@��1�ƌ��vm���/;#�H/�R�q@"�~�����t앖�	w��㵠Dw֓���]9cK��ۡ2xͭHi6U��'z�����.��bj�f"�卣1�'��TM������<��HWA-E�_���b�LI��yٜf����w��fm��گ7io�E��oX�v�/��t5��%�t��U ���������8�����U9���Ѕ�+�?� �\L-z_)
��w2��Z�9�k���U����L.=چK7�碠:&�:�	�NO2ƴ����Q5)B<�~��S^�)�#��}F�6�Ϝ䖊�����V!�����?�{��!d�ߵ�{ _/�|nJ#�>N4Ub�R�E��Wo��s��Bґ������%J׽o������N�*Bzjo[��R�9�~��!��[׫�4���-�αH��l�@"c����u�*��5#5���G� ��4Qd�t_80��*{2=T$��ku��_j�v<�� ��A�}��7�B���ۭd���澣���=P<�����*��w�	21=�j��P�h:���� �h���*�|8�'Sg숥\m�j,�H}���ܼ�u��!#Y�Y���X%A�*�@m�zߊu��gdK.(C�7�#�ߍ�Ҕ2�Ƚ�����(U,�O"Ⱦfv��ZH5���7��MOVm��U& �?/��#m�������_2��\G/��1�\S�R-�b���5�d�]�ʞd�9i��a���Α��V4�a_�ن���침č�N,��_�l�wS���2�D�%m[�}ĮߛH�#���D���n���!�ζż�ϵ�!��H��t��PӦf"�y��B7�?��?%���M���\��)�f�e�r��&46�LSa_�&Cl�t=��+?p~�����w�MFjΐ��y�S�4J�m��ʮE	�@�*������z7]����b�\�Lg�΀nf)��oqIkjM���}'%�y7�\ǗU���́�=HɄZ�	��p�dOrX�?	
�5�&M�6�8�O����<N�~rdp�#�U�z�^������+^9��QQ�p������p�X�-G�k����'����Uy��Ą�V��h~�M�kH��>�zbP���ɪp�����k'�a���=�y]~�`C$hN����GB!h����S����	��p�U�_$�}�J����FZ�%I�W��P�FoJ���'�_h	=)��1�8Cj�}�+	v�5�-�M+��-�YPh3qU���e�ϝ1��Obe�HD���J�fâH_��� `:d�����#��A�[����X��`c .���h��ټ3ʳůnL1ˍX�x�c�Ť$���]��UG:�{i��;x������T��(ӝJ�Ix�m�6MZCc y�� 9R1E��8|źp�Ys9*���i�H��P�FpK�a��1W��4���i�]B@KN��u4~=��@�_��[hIE��<��
1��M�Y�f����k98а��W(GlX��Q6�7My�`�i��M֞,����K������1�G�(Tѭy�Y������`�lq����'\f\R��Z�����p=����7��^w�Ph�v���J�C��K�n���q�h���Үa�yM�q�H���&̀\��֮�݋Z��EBZx�L /�d_�U�G�����#�34�`%r��Ao��q��{A�.��<�h����SYܿ*�t�iK���/���5ʭt�D����b�;��q\�LN���L=��*�7�t��:�q�®����A����v����~��bЛ��:IAPv��]� �<*i��bv��fv�c��x4Y�RZЂ���T���6�Յvt gzu�I�߼NJSf �-��֛la-2d�d��=��o��R$pј�*]h�vK�]�O'�p6M��c9U.7^,��VW����b�����ʬ�CWy�L��q<��>���ۚ�v��hBݝ�r&&h �Ѧ�O����~���\�R�pks�V'�/��'*9w.�"�/��%��=��]��'̓-N4X;�L���p�]%�ԣÅ���t��g�]!|B�)kh$�B�{[&kӘ��[�ۉm�5��"���g2-��e��h��Я��.��M8o��XK�A�:l:�C�-�E3�vr/Yjx�!�����y�������k�ƤR�!����vwH�ߨqz��Ŭ�.8ލ�����~����!#�ˏ�g�;��EJW���+�{j�;j��@j�7a�a#��7}#�����WPWM��ٞ32]������e�Z���_����J4���=�����{mn�=L��rYyf���91�=D�<�~<Q_�e�'���I4ٍq�᣶��:��NI��S��Ԙp~� �0LÑq���˛�Q�ym��+�Y�7��*iY�k�8���|��Od�G�_��/Tp�7���P?)�����u�,�Py�\�\��{�X��2��ێ?�������G��ɛέ`ș��64}۬�LP��r�2ǁF0^�Fq���Rv� ��6)�6�.�KZ1�>q�3��g-O�
�C���S2dM̅h��Z��Q��1��hݜ(t�Px�PCG�8H99)!C?#5�̒ЗhG���V���=����t{>��H�` ����3TU�>R��v�0��)0�Aj<+�Uh4����K�߁ȣ��ʅ����K�*��yhU�M��GP�0~*�)W�0>\��JQ����[1�F��ݱn��>=]���O'>1��z�C�dE~�Ռ6A��W���0�PK �p�#"  �"  PK  ў,J               26.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��.�E�54u1���J�{^s<I�O���h�ߪ��M:�R����Ue�wU&�c��_v[��_��6]���l	4};â.|�9ߍ�ֿk6yo��'�gx-�~\�������E#����{'��T�K�?�8�-����#��/�y����
S��|�w�����O�Sc�m�7k�1�g�����3��ᮌ�e���M�Q��4�l,(���p!�:�C��U$�A$Е�6��v�b�Ɓ߹&�g�t�5<Ѩ�������5�L\Ѽ���f�?�'��m�(�:SDvOեb@�'2|o���� x��taf��In�>���T�������e�@�Ƿ��޿ӭ;��ũB�9�f�qߞɡ�Ԟn���hI��H #�0�i�<��9i�9w̟8��:B�~5��E�*��W�޻eux�D��6����jo޶�U\�di}=i��۵�S����qM��1��<��x��DQ�����=S-n�>g��ʮ;�rC�9"ڬ��ڞ�$+�������]�3pݾ���s�������l����Rٯ�\�����٬��y!�Fj��f�璱S6��X�*� Č�o PK{I���  R  PK  ў,J               26.vec�UoQ�3m? 8+��;wwww���.�=��>@TK�EnV�~ع'��Iv$N�SJP�R�N���Y�r���De�$IT5�Q��R�ZԦ�]u�zԧiDc���=��洠%�hM���o��:��Dg�Еnt��^�$�^ro�З~�'�L��7X�P�1��d���c�Xy��D&1�)LMsb��ty3��l�0�y�O3�@o����,a)�X�
V��[-�a-�X�6���z[����6����䳋��I#�&��'�� 9�a�p�ciQ�;!���9�Y�q�z�.ɗ��U
��unp�w��w[��]�q�<����'�S�����y��[w����|�3_��7;���?�8~F���
ӢPK��+Pu     PK  ў,J               27.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��.�E�54u1��o�H�x�퓙}}z�������^��ϰ[���E��gy�=��SUp�oV}�m��՜���q��d����aQ�>̜���򠼳��P����CӏKߜZ��a���m�evVw���p`ڲ��x�%_��ϐ�f���l�&��Y��"�0�ޣ�NV�;O9���8�&�_ε�m��3��f�sb��^W��ks�E�-~�e��L�4W��(�@W|����-�Lyw�L��*��$��I-������8�.v�TN�8<�qw����M�R��>g�7sсXA2��?f̽15��$?�����M�j澽���jq@w{���Oc�{�n�#�V���^��N�/knh�j��餯"�AR'%��7�x�Z)^��	�)'��<a��|�}�\�"{�\�_�r��ߍ�wo�|8�fr~!���"�7��2�I������6W��ތ:v�q��aE���_�o��:`{��ܧ���-�1���'�D�7<-5v9���q����-�����J�L&�1f;^?}i��J�2G	�)������o�ʅ�<9�1�<�5k>����U�ƒ�O�� PK��K��  S  PK  ў,J               27.vec�e�Q�wιG�Vl�V����������n���ꏺ�2>2<�5��쁉H�"�d���-G�R��I&JȒ��4e(K9�S!I���De�P�jT�5�lԒ��C]�Q�4��s�&4��iAKZѺ0�6ID[���@G:љ.t�떤�]�AOzћ>����Lp�@}��P�1��L�1��F�c�8�3��Lbr�S��Ә�f2���an��yv��,d�Y�R���n��J}�Y�Zֱ�lt�M�c����lc;;��.v�{�\�������9��4?���Op�S��g9�y�v�K\�
W��unp3M��m�w��}�G<�y"����%�x͛�0�ڽ���|�3_�ʷ� ��~DA��4~�?�M��PK�@��v     PK  ў,J               28.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��.�E�54u1��o�p�[:g���D~�������/e�/��������>�r����|X}/����e�oݤ���g.��N��XԀ��0l����'w��2���V�Y�g�O���?�o]w���
��:f�g����F�j��_�~�#y6�Ut�H�>,Ut����h~���/������f�����nfsq�M�!y@������onl|��Vw���TW�І@W<�q���>��	!^�?$��=���wq�S��리�6���ݡ�:�΃����ݝ.���g鈙
�Q<�q�U.��'��1<�6�;C����'&��O��+���};ÿ��b�n/�|Qu���t�F��@}���40Qs���p���F֏�w�_����1�q�&M��
��g;��x��N�N�ᵭ�>1����#�~�όE]��R����Z��S��3�S�����4��:�K�VO��U��&y�F��\���;/�f���������2ko��Txf���l�G�ԝ[��N�:E��s���Cu����?u�T�7��T-�W�ܘy*��˦�>׎Nx-6飨e&C�q����fg��_�����W��?g���J^gx��*�{|qG௄k��^���QP��*j'bQ�
,�&&��01��� PK�d�2  �  PK  ў,J               28.vec�Վ��� 8��������wwww��kx >j�4�tN�>�Tw%��E���?e�Q�┠d��Rfi�P�r����$Q٬BU�Q�Ԥ����Y�zԧiDc����lFsZВV��m�&�.�h/w�#��L�ҍ�z=�4zʽ�M�ҏ�``��A���0�ag#��4/�����8�3��Lb2S��fc��ty3��l�0�y��[��P^�b���e,g+�\��[-�!���c=��&wlv�y+���v����I#�&��'�� 9�a�p�ciaO�qB>�)Ns����<�.�wI���r����&��$n�ݑ�r��<�!�x��>5�Q�s^�W��MZo�z'����g��oz��?�(~���i��OZ�PK�h?�w  �  PK  ў,J               29.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��*�E�54u1��oL8ۿM��pӥ��?�� ���3o�%��|xrc��O���)6�+M>�����������}�V,���*��}]a���P��x������r��7�g(���-������%�6>���5�!�m�Z�wڦx)�b�@�,��7��lz�B������4�M���;�?��l1�2g�'l=�'��-՜%���i8�+���4�,	t�`	t�����-�Hw�Ϡs���j��]H7l>ȸ�����g�g}�x����z7m=_�{��ٝw禭Ǣ��n]�F���v�Y�lOڡ^x|o��{S��g|�{�@�F��>mO�_6��nZ�0o��G3T��z�u�JW�`~b�N����{Q��s���ǌJ��w�?�����:�c�V//xr=e��6�U�0�\�x�����m��笽����]ݚ��W�O\�3��ǣ.��Ȫ5����+akW�lorn�x��L���SjW�&pزU�~5��i�U]�œ����D��S[M*�Օ-[V��O������%�V��\ν�(���?�����[g�1�ȾҪ�(����!h���	 PKٓvv�  P  PK  ў,J               29.vec�UoQ�3��A�!X�����������݂���Z2,2Ys���ɽɍHr"����!K1�S��:��Ҕ�,�ȣ<��$QɬL�R��Ԡ&��m֡.�ȧ>hH#{�MhJ3�ӂ�����$�$i���ўt���BW�nz������C}��D�$b�<�AfC�pF��1��Fɣ�X�1�	LdR���zS�Lc:3��,f3'��\�y�|��E,f	KY��\o���U�fkY�z6�Ilt�M�f���mlg;ٕF�N2�G��>�s���0G��8�wL>�	Nr�Ӝ�,���'ٸ _����U�q��wS�|�;���y�C��c�	Oy�s^�W���]o�w����g��5-�o���(���O~�?i�?PK*:��v     PK  ў,J               30.i��eT���ni�I	�����)�n�!���K���F@��A�C@�fx���Ɨ������{���o��s����u 	X^I�� ��;��e� ���������������@OCG��򆝑������;n^ ���0��~��\����GH@HEDD����%����:��hR�l4& :))�S ��Xh�-��:&6.>���z ::&&濪�: ���%�46���_ <��}u����'�@<��/��iX��_qp

�����WPTkji�����[XZY������{xzy}�����������_PXT�(����ohljn������?0845=3;7�����������px~��yu}s{�.4 �������:&&&����=��@�����LZ�̉��/ ��=<����_���$�s������7��X������\K B��� � ��3ȜU��T=�J���U�h!�����r�~H_ԉ�ȑ4�;�A$�é:�V1U�`����؛&'��iň&Jpޣ�k��] ����aA�9�^�zt��˘ x��QO͓i�yz�(�^�7wX���~����0���F-V1�A��K���Z����f[Yҋ�c�, �� ��n���&^]�*q1�+�w�I�e<���o�c��NrK3��B���0,#?�7�6׌�/қ�=��g�_��9��Mw�
�������k�٨+�tƭu0� ��FfV����Z�{W	�J,cG�y�����vN6�Ć]���-<�<�E!���;fA�QH�d)�(�g-�츮�~F���HxT��㬠��^%\���Mg����0���=a~�cW��d����<P��ӫ����o�a��@z)C�)֕bk���{��]ꏢh�s�CD��cT�U���1���S���wf3��h�ל�s@��D�F����0�![���3��K��C��`cLV	������ŧ/����\Sє�,�s�;��'<�s�݀���%��V.�qb�Q?��P�pi.z��8�e�Y:p"x������� FWn�V���ś]%�4<��O�X���Y<�I�o�Q��[��O�o���O ��csa���R�ˉuS�gu��Jakr�;$(��OY�*�1)��K��O���w(qЯ��Ӧ�+�C�y�d�{���\��-�G�	�uWit_܊�}C��S�O�e�$he��˻��������(@����J����E�@���o>�H'yPT����57�_�q����H��E30�_{�\d���}����9_�����t�ĭ/���F#��/���6���݅�;ժqe�Z���G!t��
�Ϗ�1cUn�~�9����R�c�;z&S�"J�0s��|v���*���Wyo�aN�ПX�)B�^I��}����y✒��5�����k:���X�׬�i�1�	ce���(X_�ļ)|���^{��o�ʣt�[rP�ܗy�'��k\E6��<��3J�[��=�L���$�y~�R�C�����&�P��u�5O]j.4c�_�X�w��uA����2�?p��z=�\�c
x^���Eϩ�- Dd
4
T^��?��7W)N�蓮A����_����P�1
_N�yh+�˼�3ց�٥1�m���uS]P�t���s_�tR~l#���&?��Ɵ_�X�߃2.�p��ۛPS�dh�_�Ƶ/��.�/�I4^؈�����O�ޔ��[0���3';���<p��x1��WV�ճI4!q�\�����������ǑepG�Ya�l8��]Z�(-b�2�y�9�h[������
�̲��s8S���
�$�~���v"��P�Quڹ:Y�=*��A�p��u.c����r��"�E֔`l1�4'nE�C"R%n'�']�Y5Ӌ�C�l�7��=�x^�f���J�F������|^v��� O����}Z��ilL��^�e�w&�pŭ���ϔ��淞���'�*J��x�iW�#���U�}���r��r���y ɑ�
 %��J�g5��P�n+6a^�Tw��*�~3g����9P�Gr��>�_��W�^�$&�43����{���,v�Go�pG�|�d�յ��{b��š�5�\+]��������5��5��Ai∋[m�H�I��n�|��?5��J].
4u��@���8�)�E�yw=n�c� ���hcqc������o2X7%�����_�}hj�&�w�ic`45�д��7���}�Q�^�@��6hBd̾޵U�|���"�������l;��	��l���H�z�
�y�/�WR�G��e"�#͡���0�'�!���	C�����):CZ2�gOZ�8v��&
kQ1<e���z1�Bn���ўS�+�5���w��Ѹ�x���ω�Z��j��I����aM6��)�(���k�m1"��Ԗl/�XC��c�ۏ<֕�z���5���۔r1�Н����Fi,�g�u�@�Z��/�Y�B���Cv��3���%,�.�F���;�/�oŴb�Д`���x$��(�1�W-"P2�R֋�O t ��W`(u�%Q�u{�KirI�}V����pq��<������ˣEw��9�׼ܻՅ�v,>�}�GX��t�����(��Pw��D�9�0d"6{i~|'.��~��+"&6p�D��o���*�Uf��k��Ҭԟ��׍bb�Kn{Aq7m�����R�w�%3�hE�M��u7GQ����x���W�O �>Ē~�\�krd N�*1�_e��ưT�=�M�?<�pt�/h�T]��``�VA[�5Nqk1%[��]�VӊR��7�7[ʢ�p}�c���&�p����)�S8�%cT�F s��Kim<�,��2Η���|�Fb������%���\JV>���dH����Pk��b}����H��:NԐ�="���#�j:��_h��=�Qg5w�����Ӏ�G�՘oE��&��{�w��g�o�����O[�4L67p�t���Cz5�ح�:�v2��cA\&K��3e�6<�h����2z�Y��m'3���ڡ��?�Q����N���mYb�W�si��N�|�=J�5Kǒ�1�c��o��v:[j��H�ɹ�;�J|Eo�|o8��ei�pp�ʎ��^54�+��wz\3̴^���+b�*<���{m[)^�-S'D+�z�;���L�{�BNcff��yF�Gf����3f���vݥ�/��|��o�rcS��4�^���+9�*�����z��~$q[��4SI����ذ/G�r��!�n����{�!��7�B�za�K���jR�Z9&1`ӂ܍*��X�1��Q�a��"���l��ê�Jչ��[�O ��7�:�m(��>��8���o�	�njL�	�o���i��c�>9��ѳ�}s�S�l�tl>jy������' 8�p�߻֬��K�,����8e���ats�+A>�P��:k���,���fc���~j:n����1�@�~d����5�@t�^�]-~wM�tK����#�e���.r<��,3������y�a�ܶ�}k+���x���zy�ya�O�S���ݨ�p�b�/�b��C�Ch}ݴ�pF:����@oZ-��V~,�SX�Ʀ`⍔j���0Uy�K��G��*�O�KsH�$��<�5`�4�1�%r�
ݬ���͟��{���w�wE�����)��#��֟��$����Y|�v���^Eq+hR�j����2��5Z>Pμ镑Ys�C_���A��Wv�'s��3��rb�8/[��M^��K[�*h1����M!�Q����X{�Sf#�
4�dX"{�"�C4SC�b?\�1�ou�0{t��iZՙS jS��8��cd~S{�j-�;p^
	)�5S�$x�����OYM���Z�M�I����z��6�x�wk�� �L"�(,�{C�r��E=�&�>���6�9r�4��|0�}���q�͈4r�,�y�TW y�I=@����YO ��� ���؆1!>��9�W6��(zt�	U���S��@��U�ޙ��6q��孰F����b�$�2/�:���`�@_�]G��8|؉]�l�
s��su�I���H��.29��tZ��M���%�n�T��QP�&��J,(�V��T1�c�R�w=|����:��2F�w��>_D�nQ{�,��vljka����*��ɥ1��`�:�i ��h�.�ù#�0������c 9"�����lQ�rV:e#��>�If��v�)ۜ��RKt1��0�Z"����'@�J��tY��n�L�H��l��^�C�!������@
��lB�sk�����S1�WD���/�I�[�8�Lߗl���?pW,m�fp�ZnG>�F�^�E�_�u�}�n*yFԘ��b�2��Pu��`�0�RZ�b/6��i�|���:���K�T*�����!m�����l�p4�ii�`m���-d��b�mX7Z��d}�f�n���q!��a0w>�;{A�RQ�ű2�s�'����bp�|bڪ���?_����!���[Q(G�?Ai��·7���sVO�W�w%��Pxk�~9����*������l%�0ɘ05��sp$���N��_$9�8�Nn��� �b�p��ô�
�e:�;�&��7�Q�[6������y�,���=,ՁR��0p?{�rբK��a����P�j�<2��y���pi��R]}�x�u�����#-�%�r	��ӳrT�3Y�M��pO ��9ݾ*ߞ����GPQ����}�u���Q>ɟ�TΈ��;ײ���Ӕ�~��A�i���]?����[��y'�B�)�������8��#:�R}w���\0�A�|�c-1���4<�:kP��lxd�d���XOQ^i���u��������݄]/ov�4�����8�`�$�Ö=������$��������X��^Q}8���~�#F��w���bJH�zA�wu�L��
lX*;�,4��Y
>=5l0��/*&����{8Vw"wOt��CiZ}�c�օ���m�ȡ0�p�������,��ѕ�liv�V��+���<K�kX��
1�MY��;���gX���If������b�I���=`�+�T6ذ�g����KƝ����}
ԋz���ȃTZ��E�Tu=�/O��?��j���i�_Rj�2ϰTs�ENe�lfU�|�n�a���)� �/(�xu�������P��,K����Y�W�J෗�tR��Q�Sg|Ӛ�AR.���,�1��
�d����
�2N2a.]$����������|��+��Xx&��K���r�9��2���W@T��FMX鼟�w��2�mv�Rw[1�1Y��F���ȡ��"�6{J�s}���q!�Y�c�zW���	g��U�7�:�kk�>?�0��p1�Ɇ�`j��	S�OFZ5�L����U�H�+�;W�}=O+Mw��B"}�ū@�t�*��6"d���"��Q�q$cE�'Gr\|�p%9��Q"�����ˑ]���s{���>h�i��S7��ip%���"�skP"D��C]IkʫS���%U����.Hp� m�¸�c�s��}�E����j�x��|���5���i������`�K2^��IɃh�������6�?�b��.i�1b���s�!�ӄ�f�Y>��8v� }�7K�:%ط6a�->q4�f����:�́�
0�����9ʲ-С��$�J���A�'�8o92:�`��x��:?��?�d.���o�J)�I#��.C�A�?Yx��{������s��cx��=Qڭ��>'�0n8�M���P4���v�?�C��b����u������ډ�����	��(����5��M��(#��/?;�����d�����S!�"�ՙ������z0���QKf�����*�3��lhN�.Z:�8o�#�q�ųê�Mm�^&˻�h�>�wK�P���'����h=�ݝ���:Br��N��c��y���e{`�~V���H��̩�x1#AQ�$�`.^#)�J�u�Xy���=���1?�UB���m�]p�w�ɉa�U����́H�R��o�Ԍ�O _݌�o��L�,�^���+E.I���;����k���Չ�}zr 1�9��gc��=���RXO�@rΒ����%�H��*l8�$��3b-�z�v	w�<�a�8r�o�;i�l�(���r2�#�P��P����e~�N�$?�!O��r�|��h'�E��A>y���%�p� օ17q��b�������g���0�<d?���|�g�.��y�[�3>�k�-�p�!Q+��x�����fi�D�}!�NW����I��t�I��Vu���q?B������;`�c8,�2�/���g��DB�_�H���aaQq�h�~�@�J9	Е4��[�Б�\z�=���
|>3
1YU�jyM�e�[2�t�\���2W���K�>|P�j|G�J���	��	��)�nU���q�9����F`�{n*�5U]��J�c[Z�"}�!엥��ߟ���\�;�1&�d�$X�ܫ���s��g�4:Q'k�-^FT
8����[+< O ����y�RFC�?��� ��A�Y��Ohc-���"T�����͖�����\��4ٲ9�UOp�Ra3U���R�Z����ט9�w�D��?�\���%���V��(�E8��[�7�$��l�����+Y_��*}|�����>9���IB��:��T/_2��#��z���"���a��m�t�W��gL�X}�c�ܿ�_�R�}Q�3U}d¡�?VD����	�1��o�?+b9�Kŵ��l3X	�:��C��N�ޭ�1��r�GbM#��HwD)�.ǵA����XQe{�)��?�y�<��g�q_���L9�c��o"K�9V���OL�qػILyA�"_dX��w�_��*{�Y�q;m9���+C.
�^Ν��V�x��~��H��������}��k�m�{�(��V������/��o}��B������c��s^��Z����<E����얰�	��Q�/�e��I̖5�g[����?���[�l	�""yW�=֑���q��Ce`6�:��}��Fo�{�S�)��_�o�%\�VRSu��H[M,����n^/�����6V�߯>���5�1VT����h�7��'��.�����$F���Cx�'〶�8Q����:NW� g\�.�;��P'*�L�K����D�q�����[��N?b!,l�r3��ޜS��A/ѽ,Œ!HU����$a{�g-���|�l��%��g�VbO|%n�Ym��n�����i1QX��3��+W/!�����:�k��>L!w'��Kp�,�B����p�&����9����^��8�6�쪸�Ѹ��3�ɕ���r�3�#V�l­�WLq�h�g���4��).��J� a���+E1C�m�\-R$��y�����=���}f@������;��%���Ĥw]�ۅ�z��f������0�����G�)���&)��'J}�:P2���mpÄ���R+g��ڼ��B�AxzN����wJ"�V�
�Q��?�I������8,�h$�޶=�a/�f��_R���J�H��r3��_�� ��_G}C�A�-��)�$�<`��
�J�O��^,�N9W�lm6�鶽_`ɠ���M�‥8�;V#��A�Q���(�|s)%�A�e[s���sS�v�R�Ma����1ʡ-\�U��'�s�,.�j���Ν��kSŃ��oĭ=�\n�Q�&3�kW���6�
J��*vŃ_��g����������WMng�;�hZ}��U�VW��#g���?=IP~=��7'�^K)*�{��ک'Z(�b|H�J��G{/Tf#tl�~�Uw5�&�R��yZ��?r���g�E��.�B�\vR-_��n�H �t{��@x�Nw=��3N+zv� ͮ�_�H����Q�����je�'�+����iHϘΥ�w���-��Ys%�v;,G1�v�ns=�Xs%��J�O��v��#g\3��j} ��^-"˒�ϳ׸����m`�"(��T�z (ke�ɧJ_~�mn{&J]CP�Z������P�������B�����Ժd�Y� �˲@�o��	?�]��'��1N���TT���WX�ŭ�35'ת���[�<�XƊ��0�}W������t%q��ع�����4UR�71���	��%�����^>K�|  #w�d�5�z��*1�~6XQ�\��� f���OG��/Q�\"��cV�II�d����2�)����
4�vUjx6I�ʊ��t��D{���(m�'_'�F���L�߷�~~Dj��yW�`��Ey���ɡ��3�������b�p����	��T�9.e�{��:Mx>���Zt���n����:��{I�i����>F�P@���r��$�5��q���y,������>���E9Dy��_h�~��U�6������ǘ�~5�R����>-�PK�I���!  �"  PK  ў,J               31.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��*�E�54u1�ï��[V���I3������_v���/��3����ߦq|�^�Q�9����Սo6^��"u��^�si]kYp����#��$�-u�������x��������������V����3��Rk�����	te���EoNӌ��ڱ������#��k;_��g�t-�����/N�|�њ8�}�!�j6���5m��󋺴:�ʮ]�����r|V�|�y�~m��-��re��Y��9=��J��~�`O���4Mh��X�4�G11OK�;�R���~g��\t�"�9��}y����Y6�G3/�[�K�t�lɾ����uvl������;�?ϩ|�r0�����YUx�ϑ����͖]+b�O�t��g�`�_�k�q풓�Q��_��k-��r��T������m]$���e�ڔI��3��|([���ۖ/niCw��<��m�I_��!�I*�n{>n;V�i�M�d{ێ�_Z�������"A:'9�/X���H�k�������j�d۬ItL�=���)v��>�i��7l��f���睒#�R,�s����_�l|��v�M�3,��o��iO-l3ԝ��& PK}��  q  PK  ў,J               31.vec�UoQ�3���!X��������ݭ�ݭ�����
ʰ�d��;'s37"ɉ����K�,�(N	J�2KS����<�H�$��f�R�<�S��Բ��Y��ԣ>hH#���lJ3�ӂ���5m��h���vr{:БNt�]��=I��ܓ^��}�G�910�$fC�pF0�Qin��}c䱌c<��$&3%��T�i�tf0�Y�fs��7_o���E,f	KY�rV��X��J^�ֲ��l`#�҈�αE��6�����b7�zI6��{��~p�C�H�;�&�8&�'9�i�p�sz�� _��\�
W���4�z7�[��w��}���x伏�'<��y�K^�ھ7������-�`~������O|s�G?��)�_��PKI�0�y  �  PK  ў,J               32.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��*�E�54u1�ïll�m�M�����������l�����|Qsn}�����[�?�3�zu��/}�����m��>��8$�5��U$ fwܚt=���c�F���3�߿�?C��oQ+K�z��ϱ�������?I�R��ԃ�N��O!�x�	~�8�����f*�����dcA���Y퓒�Oh<��~;���J�μ�'
5�|���Of\ԥ�@(hv���ܱ�c�����ە]�[e!o��$6�Z^ȓ"-ô��4_X�e,�r��X�0�G15���Y�}=��G��]��J��ګg�ؒ�N�x����9�q��kye_t��Pn�R�;����}�e٢�;����5��_	�����|�J����e79�87����Q�ĵ�d�/�"aim!)J�E�G�����"`��~�?;����{Z�+����x�����G��7d�
M�dtP��ςw_N>�h�|��͐��L�Nn�>'��Yϵ~iW#
;ʎ^`}4���m�dO�~�ܜ��JON�|�����~ƿY�&f����m$�Rٯ��o���k��g��x���)�hs��Ǜ��=�����,`VR�+b�JJٟ,�E�SW]��l휽5������ߗ'��?4�G���'�bzX$����;C��+��X�$3�č9&=��mq��CB�V��h�2kQ/Fi� ���vF���R��� PK�_6j  �  PK  ў,J               32.vec�ՎQE�}���!8�������������!<�U��TF�|X)IE��H�<�W9�P�bO)J8KR�Ҕ�,�(O�����L�R��Ԡ�M-gm�P�zԧi�Y��MhJ3�ӂ���ua�6�o���hO:҉�t��]��Ew݃���7}�K?�gy1 Eԃ��2��`d����h=���c<��$&g1�n���tf0�Y�fs�����X�"���,cy��v+�*V����c=ؘElJ�ج���mlg;��n�=v{�>�s���0G8���cv��	Nr�Ӝ�,�8ow��e�p�k\�7���n�;���y�C���x�{��g<�/y�k���s߹�{���|�3_��7�g��#
�g�'~E�PKF�i_m  �  PK  ў,J               33.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��*�E�54u1��/m,�^�U�.��S�����J���ӎ�T�w:��R�]S�3��>�e���aݚ�g��{�������+�-Wi,�ʰ�Kf^������{�����t���O~��/��nf��=���L��?�mYǻu�����M׼u�[ԥ�����ͻġ��U����<�B���.���+�gs�{��d�y�S�����ٖ�f^ԥ�@(XF�(�Nv�������l꼦]�aw��ź��J�u����v.�8��b-ϣ�@Wљ�?�h9�{�x�}�i����*=f`�_�R�>R�S��L����kc.��-2Q�v��	��k�����Xs�gwE��%�;׽�|���h���<UV�)�!��?���]B$7~�~�]�o�	�v�UZ����?�q�"����X�V�
e���/����,��ӯH�5�����4)�׳�<8�,�Vz���#[�m��qs�y�~i��^ι�>MŚSo�;�0��?���h���e�ys��վ>v-��p�u��x�e�|�����{������\��Ӳno=�~^$������
��F�^ɛ���W�(�\�ʱ��J�9X��}�<q��dRYݲ�Z���-Ix��uG��IQ��b�շe�{=y"o������o PKu��>  �  PK  ў,J               33.vec�c�\Q��w�s�m�6u�ڶm۶m۶m�H��U���L�Y��'kgO&"ˋ���w>�(Da�P4ˢ��8%(I)JS���sOyg*R��T�*ըnS�Y�ZԦu�G}�,z^#ݘ&4��iAKZ�ɢu�7�趴�=�H':�Ůk����Nzҋ���/�R^���z ���2��H�1�n���2��L`"�RAL����2���`&�����v��|��E,f	KY�r��n�^�*V����c=R��,��f���mlg;�e��n���>�s���0Gү8��1}����9�Y�ٝw�}�K\�
W��un��o��ҷ��]�q�<��c��D?��y�K^�7�/o��N����g��o�w|�?�?#�PK�귁o  �  PK  ў,J               34.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��*�E�54u1��/j̵f�U�|����ɿB�Y��N}���fֲ9����$$�}Ǿ����ְ��3�\�����M�Ϡ/�V���*��;+r�so<~+)���Ӳ�;٪_��ϰ�Z�u���E�K~����_�~����M�~�L�+�n�*�@$Е��+��C�q��}ԕ�O����O~R�Tf�1�8�@��{�&=�S:�?�q���Y�c��u	et�#3Jn��&���̈́']ѕ!��'ϙ�x6WE�B����'*1�O��+���};ÿ)o�U���XB(��3|����	�0�ڿ���^˞��zОNѩAa��^��~o���
_õ�B����\h�)��ҏ_❯�ೈ����+y����W�q<��׵}�d��sfܯlx���q�ܱ�v]k������=�����-�\&�V��|��aׂ��z��﯋;�����y�mël��=�JϬy�*g�U�꽊���_8ߦ\�&���ș��/���T��Wz�T��u�a[���.;�uQǆ_��|�\�fl(�ZĿ��ֵ7����J��rM�x����i���s��e�S�շ�?Ë���rW�w���������0���C���ZW��]���4����|#�8s�윒X[��o*��GǍ�l�< �&�!˻�s��RF�K���t;rnOu��s���L��G;�$T��^>��}C���˟�9���*�;��M PKvuTY�  �  PK  ў,J               34.vec�U�AК�v��������������ww�_�4�L��}���I&"ˋ����#��P�bϲ(a���)CY�Q�
Y.*���L�R��Ԡ�]���ԡ.��O�(e�ؾ&rS�ќ���i�'����h'���Dg�Еnzݳ=���7}(�/���b���AfC�pF02�b��hyc�x&0�ILN1Eo�<���`&�������7_^�B��%,e˝�Bo���լa-�X�6��MY~l����mlg;��n�=YA������9���+���Op�S��g9�y�z�K\�
W��unpS�y�;���y�C���'�S�����y���y���|�#������ݾG��w���PK�(��o  �  PK  ў,J               35.i��eT����C�#���4
H
8����� 0]CH���9H7�݈ "��<��u��}q����{���g�uv`~`V��J��  @��Y^xx�x������D$��$��$4�`�'��Oh��؞q0����s�r��		1r�K�	J>{!$��K@���$�$Ԥ�Ԃ��̂���td i �`����@����;qA�-�������O@HD�ϡ�!�����������g��gp�pəd�(4��Y`��Aq����]T��Gl/,\�	�=���}�����-$,"*&���9y���JZ�:�z��PK+k[;{�������O��а��O��	_��SR���
��KJ�jj����[������MM�����X���������{w�����������?\  �?��"�ǅ������.���pp���e4��a,�A��q��]��/4��,\'��	�==����߁���/���� ��K6 N4[̈́_>��(z�!V�w�4W������Aي��ҙ�e����N#�%ձ��ٻEۂ(w>Hа���J�3؂���%z�>��.��cG�0�	Wˋm�/��U6�'8	��h]����p��ӽ��Ո0�X;�ۆ[�pCۮ[�rx��@�a�B-04s��ZS��p�j��Vq*��`��1�{y���Ǻv/%J����x>�6'���'�pwn�6}���M��Jc7�C��%f[��Xl���s���h$z��-!��]�a�y�C�e_�N�o�D1�W��D����u��u3�.R+ɖbBFI{��<�@ޅ��ì�́hwH�oExN�*�{��OHMO�
G3������=����UF����7�ed}��� z�_),���|l���A��p:���%�c͠�Kؒj�W	Ll�yRSJ{1�h���ϊ�b���A"4A��9`o�8�_,����|7VWcd*/׊
���̸��tj�L���Ǖ�
�zu�Es�ҫ�!����G�tQ��ٜ[�q!u'����vKac�W�$�G�|�"�5?�S��ͺ�r}��vj�M�z����@!WJ�
�N���m�� /S��{q&t�ݺ�0�x�J+�O�b��$Q��􎎙x]�Ov��H�r>:���}6Išf"v?�1U��*�R�j�G�q��H��#��"[t\���M�.����6"~ ]�/#�G�G;�I���s��9��}�B�ݣZ*�h�*��E�Wg���Hm�����'u���B��X�|�d"7la�O�E8J^��.v���4i��-���Nʸ�Iճ�)N�-.U��ۨ�R�Q�
������u�a<���CX��
���C}�h'��u��]�H���O�Wn��@L=�~}_�`�Η�u�Ө�Ya��!� ��y9�]*�m�۳ΘI��xp�e�a�O@`ģ���{��4e�(�9��1Y�Q
>}��Z���ٷȱ�*M�W��I�1���hN����k� ��C񩚽"&8�9_��2{�5q����TWQ�UȂ���K�!��=�v�޼�P��~=i-t�Ʀq���P�1�,PWz`��~m0E[�sWT*a]�F`�A/��j��$h����ѩ�+�����k{k����SPI�)���_*`!*Ql\�A����_��5�ԫ� ��=H��[�֜���T'�x<[�������RI��|� xs��͌n�gV��`9�	|պ4ٝ�Lww��L�%5#'=�U�l�>�Itl���q�B�7I(���/��%@��B<)'�L��ƙ��s�s�����e�&̧-�Hx�"���ω���'�ֶ��y+�Ļ�5�c��.m4��kh�ь�<�NC�.�j�a��Lg[��磙*NO%	F�x��Ov(��W5��5�H�x$�($�f�K��x�Qi�2{P#(����Y�aCX����v� D�0sW=���,���Fc��������m@���A�B��i%����rQ臼���^zʢ7_��D��7�4���5>��+���ϕ����z��ݦ~�z�PS�&�5�`~V��K{�{�F�՟L��ҥ�	y�G�Γ������"�^T<s��}���,�V�K0�
A�Q*�;L䍧�U~����l��O/���T&���T�|�g�P^�%��0oQ�~i�,���JGF��u�r�����b�`;L�`��0u�NK�� �#m>U9���/�0�ϛ2��*���M�q����Ϗ���Ϗ��ȜX#ʶ�������3��1�\�U�z�L�>w=��(vF���I�'"HG
s}�a�9�(�3���Y�"�%"T)�CRc��8��6牂,���c��������j��ҽl�7qdƙ�shZ#n0�My�zTBn��BՕ>�� Æ��~L(�0���TK�
ztM�N�<�s�_�`||���J��F[x���yI��N�ǟ��S�<Z���Dл�D��IZ�(ҳ�Y�n=*��7YKi��[�}��e<sS�1(� H0�Γ6�/u��=��ϼj�v�i�9���dُ~w/�.�����.�O��7E�T�jj�LԮ��1��a��8FY�����"��3�#-Y�1k������4YDTӸ6ʛ߿̹�`�|�U��7�T�o&���UXZ-ͮ��c���&�n��������u}O[��H{c���$_k�T�J$Ul�7> ��$�.6���TÛ��VpB�o�v�iS�W@��6����������/�aF�:��G�OF������`�mɴ��ػz?y�w9�L�4��qp-g�&��>�9�&�:���n��=�܀��Z�Z]���5����G���ÇV�Ż��,o�!C(;Q��ݖ�&��?�>�_O+�ohǤk��O@◻h*I~qؕvR��T#���<�+�e��KY� ^B{g3fϷ���ѭX��J��힫�G+������V?�a�~���B$��46&]��%*�
��;܆��H�&	?�lq<7Z�-�ċY��W{3={;��ߨ���R�ɨF�����&1QC9hJ�w��2�V=`0_�/[�[R��k$������{HT)�e�N>@��ä��vI��+b�;����v�r�����T��_ܜ��aL���c&�% Qh�#y��:�h��f̛P�3��X��xA��o��W�y��?�/~&%�=W��]aE݋)�s#��WPA�v]�v�V���5sf��>��)J�t�
��0�K�����?Sus�qw"��gB��$�_��_��y�;
�ENxa��S�]*>�o(��{S�0�i3:u���d����O&�� ���R�a"q�H�}���OI?Y/F��ʸoDK#_�����ɔ�Y�Ν���6w�J�0+��c	�n=��7+�+�>�X���\���5�
��o��i�ѱa�o�?�������z}�c���^$�o��)�nXw~zL��ju5Xj�Z���(/�j��7�^Gu�:��C�����,
����H,����`�$Y��a �}U�+S�R%_�c��������sZԃ��+��"%5�x�bwj0x��Ӈl��]:,^�6B�~@	v�Ȓ}� ˌ+=�)�m�Yo<D�K�$_T��.�Vad�*\����W\���t4:1���.�e㷸�T�[�j��~�%�ƗQ\��J`���w�{�I�#>vi��y���׋�N��;T�k/�}Ft74�.6	�l#��F�w׮\�K*t���,cs,�4������>�iʑо��Ns��m�ei��N�Ӈ�P��b o=�b8X]��J�HI�gL`	(�?Z��1�0R��7a��s��	�uG����AG힐%kn�.i���f�F����Ug#=�M��y�Ѭ:� ���5�t�;���=������J��Vi��z�r����0�vn�!�тq-8-w׏Lk��4iq	^�!���@}�V��N^��k�7$
d�>P[��y&�̒�m{�;�Y��á�M�C��z���W[�W�%����i;���^5�����G⺲8֋��%�b������x�:����_��h�K��������Jȃ���<��{�jjvy6��i��5y����]�-GT�
22���*!�,�	����������G��2	O�͍G(���i��Q�irm0V�Ǩ��O�>�2�qd��ҫ����=��]��M�<�V��`�?aM}�Gp0CP������S���n=�V�VvK��F�aA��f4�T��r�=w�Rv��C'��2��& Q�%l����K���Xf:+[���Xif��P)N|�o����(�/3�j�2��@m:]�L���2tfp�ͱ��}����&K���@�G�4�� /���{h�y�f6S�6��,�zN�R�������H�}d��|>N�=L�/L��t�-$�_�$IV.ZVq<�s7<�Ќ��qY︵��ń]��
�#PuӋ�PJ>�1`�F�ك�È�c�����+K��'+$��t�0m0����[���5�$)�!~�/����j�����l�a�����;+��.�	{M����]
/�p�ﺛ⫄P��Y�u��֗�vI۾��XR���ßߋ�,�+��Ѓg�{��"�k̄1�l���r�%�+�����_R[K	o]{�X*�����+�f��=ygȆ��|��q��Os��'V����s]��D�Xg2CƿP�Y�:��|����|Q��w]:�n���}B�����u��CQu�,uB34��r帢��9�6�0����#5>���(���uj���k�E�ځ�CB-t��b�3���X��|*��{��B"'k?}ŒC&:�$��=B�!x���;ڝw/��FA��u�(�8��|���x�6���ȷ<��ne����װ��n1�>�_ۋֽ�����(�
��6�^�4.���iE�a�q�-ۦY�q)���Ηz�卼T�vĂ3��j�mތ�_nE�8��kp���	�~�2n7�Q6v�IA�O�S��
����g}����z� ���5)��y��=������O�
'c�H�J��9�d��g� -�ڄ������>T��;o�\��$8	�Z��As?������W�m���Ѯ�>��_�k��솫�����Rc�;���M3"�)�q4Ĩ�Au�T���&6�������=O��?�Gj�FsjB�8�,c'�����������/�x����v�����Co�?�jD��3Yje���r\a���rF~�)<��bO�c��KyB�)L���9ȝ�� bX�2!�@{e�E�K�r���^w��uET1C�=d #s��N��jk��!�ԁ{\%Ð�(����μ��V���[�?d�\�q! ��ʣ��W}�[�@��&շ���C��>C�HE:��G8��кS�Ac<��P;秿W{���˪����^��x��O ~)H�ػd���A�#;z冶N���|�:�:���"�(����5yhVK�- �'�~g��ZƒVgѼ����o�u������iE�y�.q-��$�K7�AѓE*��ۦ{�c�Uj��
X�:R���X�����D<�i��p�4�?�3�٦3.�y:b �Xj_��-dG���E5������sl�vN�gE�5c_#�lv	<WB�kt@+�>��P�xQ���\�m��Z�~p�͵����yt���2-,���6$~��2|VP']o�O����[����"u�����,P}���4&z����<\4����3`i�|�g�T�H�;�%,��y��^��ǂ�S�_<[ˮ[��?��b�Z�����w�G�{��{Z?��T�p]'�GPIt򊖹�8�2��Cs�@�i㸯�+��q��L�$
!D6�bJ�p�9�����܊o'Cn��y����>� ����[haͥ�e���]��Q��	=|fv3U��#������z��m�Q�M��<[�Q�k�6��Wu����X�>(��7D3�<�R�gSC^F�v\S�8�(&��LT�6��-���z/S�d�}�K����ͣ�-�tT?�16G���D�1��|�z-L��\��՘4
>��6F�fC2�q8	~��SN	�zc�㬬�ў�˳�JS��	�C7��3�%K�/Ex2�9{ՠ&�"�����D��z10p&uۘ����5u�Tw,^B�� �k��v�%=�\�K��<��!=.�`�C��[#Y�5	��v��\�����z�R��nm���{L!�ȹE�&���%���K��l�q���P��o�S���04s��k�����6�:������wT02ai曷-�}����Q���-~�]��p�ԟ%�s�$B�8P㥝[�a����q�5WA�]��mզ�'R�|�%E��ΑX(%����c� Hjt��d�0����U2*�nsP�LoE�rW3v�n��}N��Aj*��0�77Ki㚕V���0	9���*F�@Z^b &;~�d�fe�V"�D��}�R��#�n�Rc�sU�An�	�'h{�,1�� �؋T)�{<�4?X����^���(�y{]G��zj��"����+�b�C�w�ϵj�\�JO�6��igwןi���Fd�(�����n"M�y|r,=�E�3�����?��3i���pp�!Ht���0�C鶵�>��%���1���&]�u�q�WZ7!ZRlQ!b?���X���f��7;*����D}˳���hޞ}�_o�%�n�i��:�
��(.�ϋ3��$��.�1Xh��2��2$��l${p���qyvmK~u�g�Pj�bn<뼷���l���)�����n�xI��V*���<,�X����rN�ޤ�!ewf�f��_� 5�J��4mR����b��<���O�/k:R��s�\�JAQ:^?67��ۿ�$9��'�a=U,7?�ߔUJX�A��>g	����kO�Y�:��O."k�v<+/t���?Cg~�����p��o�s�.����G���VW�7�0�\ͤ��&��mZ��bӋ�����'���0�N�*��d.RV�/�;iS�J�F���)����r�R�ЁD&�(��8���3����λ���UkW V��� �r+lm�bS=��1	m�t7�	����hv���?��O'���9�韈E�
�˲�6��Ǌ������1@��$�֟�x�R����9�^u<��܋�$�y���C��x��T�p�u]\Iޮ~Pvm�1�Ѝ2o�gza���L1
v�����#/+��v)��:������ś�x^&���_�����ŭ��K�㓥)|3�� OkSoT
J{��U�m�狽:-�����{؇��
�a�Bm��:1����%����#��4�$��7q̓��ТR�I��H(�D��K~�v�����s��ӄ	��x�F섴�-�P��s�,ߩ?y1�kG��vTO@�^0����>6[�"e�A�:����h'�T�u����b�
�aITS�T�B���y�S�ܮ��I^���j�{���2�`��8�9'-�<��B��H� �1��<cG0\����;��H��3��Sy&$��y�8?�1\T\B��z_�����R$ޜ�.D���	�N����u�$�lx��{H.�5h�9ž��_`�Mc��X�K��������C:ڳXO��z��]t�y�b ����vo���eXy^cg�)�}��9R9�̲��'��\^�Z�Xyu�ꪫ=��߾ڋ�žr�\��b��cm�7B�W�e�_��1����o��.��1VKcD�⧻O�>s֊�N�ج٪�B7�u��5x������@7Z��:AM�OU���c)�˾�I:ׯ����H��z�h� J�v_�,`��E��r�Us)ؙ9�=�Ҙ��*��
Y�#vQnɪ���GQ�xr��VBe�T;|Tp�5ޠvV����;A���e�y�w���T�z���'oH`�ˏͷχ:�q�淡�������A&�R׌Sɲ��L��0}�F�s��+4�������dc�U:�<[���Q���G�DR�uD����/C�,�(��7]�7	��n"����x����MN��">t��w�^��d������mO&��?�2&�H���2�{��ۤ_{s� u�,��u�P#/���U�����Q������8�f�z!�WЮ���9����ɂ�������lf,6~�=C�4F�E\'BM�e?C0�P�\����h������:#AE��UƘ@D<OFe�Q`������!�"G�s�{�-��Nh�u�EVp�sr��t����Ę�y! c_dj���Ԟɉ��~�_H>䓣�ȱ/�zt���u�C_��2�v��-�Bg��a��ع�Ly�u�z6�Y�j����6���q7gU�
���D"��G���6�1Nh�I��q���|�+�а�c|���ٜ�L&�]�}|pDI�G+O��B�[r����5�����1�S�a���6~g{�Q|*L>S��c�{��DP(�}�ԇ�F��g�g����Kq/���"��\��d����Tj�}ʜ���r��:�Ю8���K :��Ư��!���zg�m�k�_���i�y���9	Xm4�����"����L�!���~̤��w��x��Ѻ���\X`���J?$r̷�X�X��G�%�5/ː�%%J;���4�%��J���|d<3!!����9�+�����`��o޼��z�����D��S��ٗ��*��)�-��tZ���F$�c�PK�3\�l"  �"  PK  ў,J               36.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��*�E]E�`���KSv_v�X^����ڈ���6|���f��]3L���5��/������m��P���[��zA��3ui'��:����y7G���4������a垬��tm��9&>?��Z~���܃k����f���Z��a�5�(��CĘ.t��CM}���>�o5�IT��e	�pl��Z�&	�wXʟ�t��7׉Z|E�����8��h�#����3���z��u�k�
�P��i7^x57�\[r��ڄ�kV��:mx"Hڒ��kw�;�.,�SXԥ�@g̔=�f��"3��,%�O�_Ʈ�|ȹ&���w�x��y��{K��ko��)h���kҩ[-뎊nl}���ڲm��ʙ�"%4�������*�9�����6/��,�\tDᗀ㿩�I�NY��cӴ����yr=�����.��d�r��y�>�\�wE�9%o�&�k�J�c0w��w��͞�;�ߨ��[e���l��-�M6���`_�4��s�ͧU�=��ڽ��hzm���S���0ٿ�T�u����S�x��n�Ɍ�>���w���/��3\p����2Oi�v�U�6��U���_����'n�/���U��)�Wa7U��+�`o:��a�C�Q7ϕ
1�9O���8�k��;2��$q��=�zu�s�M�M3#n��?��ː�dJN��Ø�=��N�\���㺴�ǌ��9�^��I4
����	 PK�.
�  �  PK  ў,J               36.vec�ծAК{8@p�����������!��k|�4�tV�~ة�tDV����Q�<E)FqJdY�4KQ�2���@�,���T�*ըNjR˞�f�R��4�!�h��h��TnFsZВV��m�h��h/w�#��L�ҍ�����)��7}�K?�3��� ��`yC�pF0�Q�N��7V�x&0�ILf
SS>��M�g0�Y�fs��|�z�E,f	KY�rV�RoU�Z^�Zֱ�ld�SĖ,[�mlg;��n��7��}z����9�Q�q<��z'�S��g9�y.p�;_һ,_�*׸�nr��:w̻��>x�#�Į��������y�[�齷���O|�_��w~�����W*�ߑ�PK����l  �  PK  ў,J               37.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��*�E]E�`�w�y�6�G�E�d�yu�̜�i���3��Pv��� �\��~e������n���������(,��`����^6�f��]�������V�I��N�����M�d��2�L�*-�ۡ>��G���r�k<���fm��f�.��."����߆�S;~_�x����7y&F-�4l��t���ܝ�V��:��<a�6U�U^���z��2�5�-�Kc�
G�3��7f^x�#���i�tAd�x�FI�k��*�����{)��?���[[�&8��f8ѬX��ֺ.��yr��E]���g�.��ԦQ_�^~i�����w�s��?%z,����3�'�?�X��xl�ڪ'.Wuiyke�<�b<�Y�}�[���͇o�Q�Lw�������뫗��F{�y�WB{�\#�Yz�_�d�ٵ}#�bu�~n�̋��?���6�j�Q�-��%�I�j>�N���m]*]t��J�������Wf�?>�puof���#��k�9����g���e;�7�q��P�{��o�f��>����P81r�i1�g�s�75;�dֱ�O�\{[Z&��;�������a[��ք<n�.]��H�-m����<~���o3.���#��x�埠s�Y�Ƃ�),)"�Gv��N���V=�I�-3߮�MTo���G�YORc���u���	 PKY:�_  �  PK  ў,J               37.vec�ծ�P��{8@p�����������!��k�S�f3H3�����n�D���Q�<E)FqJdY�4KQ�2���@�,���T�*ըNjR˞�f�R��4�!�h��h�LM�f4�-iEk�ж0�vY��r:҉�t�+��n_��r/zӇ���?�
b����0�ag#�蔋1zc�q�g��d�05�c��ty3��l�0�y��[��P^�b���e,g+�Ve��5�e���F6�9El�/�����v����ao*�}Y>��8�!s���x�'�Nʧ8��r��\��|I�|��\�:7��-n��1�r��<�!�x�g{�<��󂗼�5ox�;�|o��#��������?#�/{�"�PKu���p  �  PK  ў,J               38.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��*�E]E�`�{R�~]�_�;������Սo�J<��9�E0{�y�wf�����f�����6���sT$0�CcQ>|g�T��Ϙ����?��pm埔�Ϸ(�^��a�5q���u�Jj��E�>b�|���W}�_�N]�$m����#���W9��y\UB��˕zO�e71Oh<����W��İz�}��q�5�5M�E3ϩ���[}�J&ui�ta�#���hP^ha�03]�$G�LC�D��*}<m�}��ڡU�muqv�w����m�x2̚O�<^�r�)�f�U��|��V��o؅[q�N7�B�,Y��VU]s���Ea���{�f}�q����+bp��y��^J�9�P5_+�EKM���ö��W����Iai����J-�Mc�ʍy|=���Y�}�,i�"����~m��#z=]EB��.'�y�ܹ�+��3�z��oA�ś	����l���Sۨ2��JI����������Ӹ�+�����DL��w�\.*��{�v�1�m�9�V�R'Ur�0/��A�ں�;�_|�&ɖ�4��b�'�V�3O=~����G���-Yq�&F�|/!��~�?M!���/MR��7�۴qQ�O�፲������ʛ�Xr�r�Y��4򚀑 �t���2�gRk�n��}����u~���ז��7�
�(>�sB�>?����7��T��� PK_K��b  �  PK  ў,J               38.vec�U�AК���������������Cpw��O��9dr���Mu:��E���ϧ�E(J1�gY�0KR�Ҕ�,�(O�,?*���L�R��Ԡ�=���ԡ.��OҨ0��zM�4�9-hI+Z�F�m���ܞt���BW�����C�I/zӇ���?R~t� y0C�0�3���J1Zo�<�q�g��d��\L՛&Og3��l�0�y)b��y!�X�����p��,b���5�e���F6ٷ�[l������`'��͞�7�f��'�� 9�a�p�c�O�;!���9�Y�q�)��z���\�*׸�nrK�y����>x�#��x��T~�s^�W��o���{���g��o|w��⧽��ߑ�PK�$p  �  PK  ў,J               39.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��,�E,��`����=�WF��5�U��~r؞�3������p!K�[n���]��C�/-����7���R���V�%�5��U$ f�{�խƩ��-�n��ӯ7�v�����nB��&�+=o]�_N����鑵8{S_��S�&�%]t]�*���b�z�{[��k��К�L�~�b��e�w��'���u�����������^���y wsi�Ƽ.�e�>��7f~{cj��I�d����9����ؽ�eӦ�0ݮ���/�ԝ����6�ۺھ[:��,������iO7ui,	ta�3f\�6�;���)�Bf~2�(��s��߹닼��沇�;�,���m��c��ߧ<n�y4(�U�$��3U����'_N~�8��ڗ��tyt<X��{�������'8
�_��#���;ۂ��k��\��:X�\h��X�v��E�����_~_/��=3�D����_��#���P�����>w����U��x�.n�ݶ�Kjo��M�f����xk�r����_��Μ(�y��1��w����>�S�.Y�JA��}����f���v���se_�YUM��{�>�;���ˮ�8�^(��%����h���mּ�f���jn�%|����.s'`��2ui,�]=C�-��1�?|�,�++�쿶[�U���)�KZ^�E+������ۥ$����M PK��?^  �  PK  ў,J               39.vec�U�QF�S3�@p�����������!��k�`rY����/U��,/2������E)F�,�nIJQ�2��婐�GE���BU�Q����Znm�P�zԧiT�Ec�&�)�hNZҊִ�k��h��Ӂ�t�3]�J����z���7}�K?�3 ��@��3��c8#ɨT���豌c<��$&3%�b��4=��d���\��ͷ[����,a)�X�
�]�E�ҫY�Zֱ�ldS�؜���mlg;��n��?��n���r���(��g�8�Or�Ӝ�,�8υ��E�K�2W��5�s��ܲ����.����ǩ0��=��x�^�׼�m�����|����W���7��?=���;�?PK�fU�n  �  PK  ў,J               40.i��eTP��g$������B���nIa�i��nA�����^�w��r?�{��x�:���;��O�O��W�P |  ��i �@G��a�@ LL,l"�/��	�^���^SR�0p0�б�SR�`a�����3�
r�p��r�� &&&�Kl22nZJZ��g{� �c �Y(@:�| 
>� ~�'��?������١���*
*����= ���K�P��Α��/&�^���X��	���?&	)�kF&�7,��|��B�R>B�e`��j��Z�:�&�f��V�._]��=<�������'$&�HN�����_PXT\]󫶮����wW���޾���ɩ�ٹ�k��[�;�{�g��W�7�w��P�����\��\/PQQPA���p��>*-:��2�#!��dLvU'&=��	���_,����A�o��;0��/�������(���� ��Pͭ��@�ߩN\��	�G�J�dB�����2����9\	F'�$u'GU�? ˲�h�O8�-F[ü.D�Y �y��x�_�[DA��C�LKlc7��?w�=^F{ށw�x:�I��M�}o�g��M���K��c�^������D��C�j�v�]�-��'f�"w�QA�菽MU�)^�
;�e�Ή�IO����*)�x��K8�2���Mu�8�c�>�ٽz�����+�/ȣ�����X��|�S�v9���	�K2@��pf� 4��{p��(�tE��!#����i��ok�rP��9���@.Xk�#�ōO�1+�%����	��yb^C����p�=P�x��jO��)3���HB�� ,���Ѝt>�˸�yJ�7�T�h��Oq)1s����E5��3���Qb
b�
���z��T3'���E��!bk[X|�Cmͱ��"� :�
*�G*��
�.s/�Rs"�V1�ίЅ�h;:z�"|�[������l:0|6���u�uEg�37]|ǥ�&�z�Q���U�U���&&���.���&�W��_SC'���Iv �Ή��#3�O"��>hԍ�,ӆ>k�x�������O���)s%�@	.|�KS �2g�K����z߃�t�㋘NE�f�o�|�*�-�I� s��K&Z���3HkM�x=)Ç1��[K:���A�'�/H��Ѱ�{<� �I7�##�We�a4�u�sռ�y�L[��R�ͥ���:���z�3E�O�je��P�|��щ&�6�(��/�8��a��"�P�,̹��U5A�e�u���ַ��{opC��$L��dE�4�Qg����9^������X�����i	$��qFl���O�l�X�� {+K�@^�5�"q%��=p˿Z�=�������w����5�fWY����iz˼g�E�M�����V�5�~�(gZp�M�	7�<-�tk�m&�12�`P��*dL7u�{s�F��A�`�r����rN��|8]����Uf�1�;4R$�*�v�ՠb�J�-��;�e��#+��p����:���lX��_8U'������Tj8�uPjD^Wn���; �y�R_�MG�m�M~i�R��@�bN��z�\���A�a)�d����b9ڈ�����Zৼ4�@KukR�Ic'�A·��{nG�($6���X[�8F8]Q�����0���kE��&�,G*�e��i�e��W�E�D��&&�l��,a(O���<ڍx��t�|�y�S2l�'��l�D���_�Ʈ|H�����j���'?�1���p:xM �i���M���FdJ���{B������� �� �{uL���Q��X��ó���rU�Hn�m��lo�o�_��\�υ�a��*��̾!��D�U�پ��1��֠��Z|���lg��]bS4SX�Ge;N%��T(�J�8��c��>P�}�
D��\����zW����UX��l+N�H�������v���S��IqX���[)=]�$�����M\�~A��g���cx*nK�Q���XQ��t����C�t,D��=�( Ɯ�v+aN�~Li��1.-�+�t�J�j{�뼙����G���`�l�ܭ�}W�>!Z�>?;"���Gk��� ��i��jq��c����6�\��y�T��&.8	�J�ú�⬡>��܏�|2�%q��E�!��H���"���_���/�a��
}�3'S�̰���(�%�[�?�J��Īy�pV�t�	1->	�	T�dM���� �6�#!�o7X�F^�L�L@�s,��L[,3�
�%2���rן������Fq�f@/�3��Ri���� T@�gH�c�|��	�V�^�����[��ܷ���A��Lf���h��{��k�����Sl��E��{�����Y���v��t{F�\�k���Ս��OQ�)Y����#��)/Mb'����`���`�m.�X�JV�ׁ�s�0w�w��48k����;��.W�ل�H��\����"�rO�f�]GI��;=e�UE&g���<R�g�K���V��,������ U �Xk�����˪�0t�E%�S~"�paSzȿ��<)��yuXv1@��ﯶ���8��� A���[�_~9z򆨶�2�ҩ'�U�y�ʀ�_]beГ�2�~�e�l�o�?z���� �9H�P�%Q���N�x������K��PV<5Α{�1��G��\�N��V#�So�nx%(��r�/`��֜pئ���"� *�}J��p���-(�8F��EI��}y�	�U�����ȩ>����Z�aQ�5��shyk4�т��ڧ�$@Q��Ҙ����_��{��B].��i�7�Y�@�� 6�������Dmm�{/*}QZ�4?;P�h�e�r;5�����7$Gޅ1yU�š��+��8Ӄ'%�_��t�U�̧0�O��1�_06�|j����	����_:�Mg%�j_�;O^��D�f�ܒ�^Y_W���**�~��;ݷ��]P��U�r�RЬ&faM����6�ݐ�B.������ݙ����Yb���M?�
�2A��2G���I
�-����F���ٓ�tbQ��^��7�c��%\Uh;�6�O�i�>��[�k����ù��s����٫*�?�OcQbz'�zu-�t~0��'��Hʮ)I֣�H����4=}��e����]|Tז�D	MO?a��c��gY�f���:�����}�#��׽�I�5�p[�UM���xllkX2�4�ǨUm� ֞ܖ��n(g���'@�G{���[6j��q=,M��t�*F��< �^�;uo����I=Z�^��.� �X+�~ʆ=� �"�Т�&Z��f	��M�@K�y9�҄)�+�?"���ys_ii�N��=y�q����5�Nj.[f��%sF��Lb�R��`Yģ�r~��TWg�F'\Y�Je�v���7�Kc�G���ɟlq��!���G���{)��l��1���;�g��=�}�E�/�X:���η�!vSFER,����P�%_���R��vĖ���I���--��.�y�4�M\���h/���4��)I�L$�`�}����1O�}xWg�W�oa�������b���i*e@:i���x��Nk��C}�G<�՟�b	�+)��M�F��s"ۅzk�^��PC]��ΫC���lV�d��=\�����y�!�iSﾏ@���IZ;l/jJ�%?�0��KDp�-nGΖE���D<��O�W���
5v�3�I$�%4Yt��e�ЪvW.J��ÿ�T8L�{݅đΕوw��Qu�\P���}���;|�k��=�s�{����D�X���kka������3��t���F�5y�E��<j@���*{b�0�%� s��X8��ןd]��4�Fj���,О���@�:[eﵗ���dsb�
��5=_
����{�b�m,��u
������̔?���U���� ����U_�3<�%���H͜�rm��st�Q׎�hH�c��_� �����t-Wg>��,��S_��Hn�[cڹx�_.���K@�K� M��$-	����9ks������Έ�8lFBGV�'��f�l9��X�N����m�ff�>�������� �%?*��:�����6�vM�M�������|F��\)��()j+�)�,(�,�O�1%�$l;�zg��M5,1��Z���K�[��O@y����(x����4��Ľ*���F�����D��t���'�0����@NJ���|�sr�?�"�c�
���m���2k�[$��[ޜ�����u���_�E,y-�x�;��(Z��Ћr��FF��`��kڴ�ֺI���G� ���ҋ�4S��
�&8����%�,���${n�ؤ(��i^�B�z�T5�q�ITQ��V��ǌ��Ay~GiJ�N3���X��;��V�f��3�n�g���S��Q�c�3�!W�$������*�P�`�����M�e�\�&V�b's �L���ӣ��ȷ��h�Se����-���Ը��_F<���}"�3v��s-'|����nЛgXM_t$\�V�\������Gўt^�I��87�aѝ�����To M�i᝕��pr����.����^�����2)�Z���]�M� 䫁�+�a���zÅ+��B�Z\eu�����G��a�ȏ.B/'RG�K��߱��]��-�g�!��H��Ј��s_����8ňt�P��W�ʌf~�qd+�(�|�����U-3�"���y���k��B#L���Mf?c�3�+���0��
�kF"O��ۄJ�9,�6�<A���^�Ա���е�|o���&�S$�+9����XɜޟI���3:㍢E��, �-Xbbr��?�@��ҿ4^�3��J�����ɽb7ݣC����1��;�y�Ot>v=۶-��P��Ʌ����N��`kS|0�?�zq��z��[kҽ��f0!�����7�����zWi$h������\��+��/��d���ZHZ46v��vV�������̈́�X#3C�V�v���aS�ݠ$�ј�E�~4[�)}U�@D�Q�z��
��9�X�q���M�h>�A�^��b����xl���܄�����@&���r���&�c�|�r��C��Yc�r^�VK��~\�M	y��"a_Ce��]��]�H~AK$�)�t$�]���K��2���0u���c�vh�k����c�Fn*�5#��p�O�E�Ѯy��/j�˨2�S�G�2���\�biX�� #�;R|qjh4�T˸H���&ŏo�W��� Q�me�y�)�&����^��]}�?c`m8s��ѹl���|��Ż����0�T�߾�#Dx�z߯��+��6�!Hu�&�����T'dQ�7"M��&�Ǫ2E6Re���œ�2H��*�t�ቸ��'@�5G�}�9^|�����ew��)ަ�2c$��a���S�Hq�M�.�f�-��]5|}���./S��On��h_? Dʔ=@��i���?��J�J���"2mN,�i�Z9aȢy���V��k�LǘG^�' �r���8գ�#��x��'���"����k[DJ���T$P4�<��V�	T�\��z8k�"�|$� Y�#�vFLD��]L�T�j󸤏�@�-	�<k�<��'A��2����O�͛�fa���C�2�
��Gӗ/�ͣ��.\�]�cr%qا�Ǌ���o��5��xI	��59�Δ�F!�cB-d�V���{��AFCKW��(�	���Ea!�Fס���],O�~�������m1?+[���<L���]{>���� ��x�	�/��I���͆1�N�!.3#���խ}
��l��VB��|�n�t��ygoqRbr��7�(�����0G��������U���M�-��	p0�H�*����|�0��ld�d���
?e�՗7������7�*a6�#��H�R�j����1�f+����tfs��E�|��.!e�'*�]�����d K=η>��[pns�1��'j=��z��=KN��0ښ�)�p�v��=)���{C�W5�KQ��țaE�p7�h�����zY
[Q� 4�P�!�!,��rD��yH����?L%�&�����!ӨE2pt�3 {u���5u����ߣ�S1��]Γ��困��!'!��� Q�M�N���HD(W��f���
����Z5�Rԅ%ҙP�FFx~[�Ք�����_�y!T��E��q|Y�C��Z���J�v����5JKF��8��I]֢���*U
{~�/�A� u�6U~�`������+�)���?�����\�g�f�̐�i���O�t{ �6��q̆XQ&F��-r0��ӷ#�NeG�u�c0������U
�	���eM�4�L�8�4�tT���r������;�B���!_S�zX�Q��<���&��ͳ���P�:x�����I h�{|epF� �{ �j���a���QMCW�R_7N�����D���X����
B�,H1z��_��N��/Н v���`�<o������y���sֶ�c�l���G��=?���u�dԾ��H�F�kkwS7����x\���b:,�`]�Ω8���pv j$I�s1�`k��'m���L�2s50����#���~'�[�>�6ݖ�FCN�ڃ���[k�bt���4�<��\O�_C��ѡ�D��d1����S���3����h�(�VnIN
Pw���Z�<�
"�ތ��Ee�O �,@�4j�b_[�!��O}�Fx��P����-Z{����[e�m�TT/���]6�� lf� �iFi�D}��+�-�z�jɡ.m|�/��\��ڱ�!�L��;��JK�cs�;*�0��^@�9�T��_���X�l��RI��ykc�M���l�.o�&Q"�T��2Ś3[�VX�����%d��RM�)�N�����fj'�t|�`HY�� ��2-��'��Fx�r�-��K�Q;�EM-Y'�x�R˘�d���rc��J\�m�Q��ZןL�����j	7�IblG�yp���Ǻr�9eW�g(��@'L�(p�p��O!+��(�ܴb�^֨�����`�N}H�]�a޵@��Q=��=������_~�bn�����a�:���3��m{��5�n�iq�J�� ���OZ�\���A�]�����#�K
���v�0��cO�"�譚�b���?ב�?KxbY���,�(����64DW�vB��d�˻܁�V	fT�}��/_o����UN7��׼9YU�D�ӭ��
�򬮂���jH�B�F~���Q/>��2y���<�qG���j�<ھ}^���q@%5�ʄ7V���g��ө:q��5��_ώ���εŜ�Q���d��\ǌ;��)}�`�v�Vf��N����	�!ސ`�oӽ�Vͅ�,�7��d�7"|>v<8}H{����]���tQ���!Q"C�X|e]�ȹ�H�Aذ��{_�h������5	>�S'2,��CH���U��7�#�y B��>�.�g���1�� DS�:6�40ܱ��XI�.�	��[�Z;z}�+1Sq:������8u��c|3&�`���H�^J�Go6��L�����b�'��9%x������!p�G�q����f�4��v !~�v,����7�M��jt*+<�����)���z޷��}�iP) �+��zB��Зx�#���+d�:졤+~�39?z�! �V���s*}To����xn��o(9�Z!̋����=�V�����XC/<-�@
�#���U&v���1WBi>H�C���M�}vV�v��8^5*��Z�m��0�R��?��������_r;� �; �6	 �`��MqŰ6�^�@�P7����q	}E�� �浾��#V!M�~1�[��MO@s[��fh�G"%-M���??9�;H��*�c{;P>��t�7|�v=�{3a�.�6U�4�0<f��R��G�9���[\C�s���V���\���܇P�;��|X
z�Up�h
�@u|`��~��$O"�o��*�RfQ}�fRM�F�q���@�k���mms&��?�(&#��ٳ�T�ԑ��n��)Oj^�S�����o����IZ?>�v��O3�� �o���LB������/���T<�JV,��ɡ��X�cl�ߓ����|��  =�W/���L��%}\"�۽\9�,,$~����hB�%�U�k���68�-��_���'s���r*�S�^\'%'8�ʻ��K�ݛ�����1�,���>�&d�Ġ��׃��*ѕ�oɦyW_>�����*-(4�G��*��?�v�~�������E���K�U�P� Ĳ���j��r�J�;��w�0� 彎'�/��/X���#L�~Yl�a��G
�L[2�"n|��,G�m9&�ǫܫK�|�}�5�N�ɹ��)e_ .���R�|Ձ�n���i���_D�sҾN�0l�LtY����[�-��m�a����E{��ӡ�����<6i�y�����k�l�>vT�Z ��#yHMd����	H�|��Ȑ�����{fG;���������E�[�I�����⁝�eᘜK/�X`*��!tE|���p��~Tv�Ð����A���t�e�fj��%_��������Q7|RԗV+6��T]�S��_<{��n
.#�N����Z߸��׏ʳ�WK0�ɳ�HN���aJ�k5���/PK�(���"  4#  PK  ў,J               41.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��,�E�54u1���6�^���������0������3��*r<mG�qA������3S8�f+���[�ɚ�3���+XE�a��2��������X�禮����nf�It9�dX`?q�nP���P�w��G]ת�\ԥu���������<#ç?O�hʚ�����G��
�_7��r�G���	G&��_�Z��Wn���!�¢.�Q<�1�ź�>�+N�<�7g��lߧ�{�"���bni7C~mqxs�폍�j����U����*�Hg�����mMo�߂���Ow��A���-���b��ǘį��]*}j?��dj�����P���W��4����L	te�ak��kK�����_���3E��f���'S�	�.z����Y����O������������Tm�\�*��_W(W�Y��I��6�}�5K:�NK���b����0;��P��&o�?W�,;|��y�Q�?Jm/�4-� y�o��K�[�T⪞��{=~"ox> {��E���=��1�Xg��m��'��7PK�T�t�  3  PK  ў,J               41.vec���Q����E�\˵l۶m۶m۵l�[�S�t�g������=Y�9�G>(H!
�q��)AIJQ�2YN�u��<�H%*S����NjR��ԡ.��dQ?K�@7��iBS�ќv-�Z�ִ�-�hO:�)�D�,���J7�Ӄ���7}Rn��}�t0�AfC��b��=�Q�fc�x&���h7IOf
S��tf0�Yv�����c>X�"�$e��;���`%�X�ֲ.E���c���&6���lc;;үؙ��.��=�e�9�A�v�}�c�'9�i����v��y.p�K\�
W��ם7��-ns����~���P?�1Ox�3���w��{���w����go�)��-����7?��H� PK/�&s     PK  ў,J               42.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��,�E�54u1�����mYa��������u������w�_�1;�m����?þ�!�L���;���n�>�f�.�E[ui��L����n�K���ζ�&�_���1��3���-��8g^�\�r�����N��t��[��]}Br��HhC��̸�X�[�P�[H���^��MrjrcX�����?�!RB�-Va��b-�bQ�H�+�(��a{6�mY�~���fݝ�Fr��⃑i�\��
����$��_��]ɼ4*��լ)�����"�t�lsOޛ,q���c����z�z��}�z����o|�O���a�B���jkD��M��q��M�_�1���,�I�>�u9^r榴.1u	�2�yW�_r����r���+�EK ePƒg7�ݱ`�%q��yI��'Mg���`�}���������N��:���}6��V[������� ��:ۓi�֬g�*�}���V�Y�2���?�L�����<��ʶ���Ҳ;bw�>�0�3���e��Ev��j�Qj{Q*�˻kM4W����K�Y�1?�_��Z��-۵��6*4�c�R�޳G��R,�����	 PK"�{�  M  PK  ў,J               42.vec�e�PA�s_�؊������������n���� �SƸ���6���,'2��.y�S���h�E1�8%(I)JS������Y��T�2U�J5��SìI-jS��ԣ>�d�0K�HnL�Ҍ洠%��Z뵑�Ҏ�t�#��L��]��nrwzГ^Л>�M������� 3��cxʋz#�Q�fc�x&01��$����2���`&���7Go�<��,`!�X����e�\^�JV��5�e��6d��Q��f���mlg;ӯؕ��ny{��~p�C�;b�Q��9�INq�3�MY��;/_�"����r���zü�-ns����>�zh�#�1O�Χ�3�󂗼J����-�x�>��|�_����wo��3�?PK0o�r  �  PK  ў,J               43.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��,�E�54u1���;y��<���`O��ؚ�;u�N�����f���,ל����|��V����n����R�L?.�n�*�@$Е���|�S��k������?k�{]���5K[�Yθ�J�O\]~IRq�SQ2��_���4Μ��*�K��o���ip0Ӊ�_aN�k����g(+����b�ՙ��j���ϑ���wt�ƢFBf��QL,U.���M2�[�&f����v�<��FW G��v���Ey��8�)�������W7�lH��'y����1'�]���?��SſO(&O��yr\�c���g�e�3��i<]���4�=�gU�W-�c3���Px0q�/}���woz��;Qz����]!�b>��__��5�I������لKcQ���g��=/�i�7�+)a)��՟�ޟP�4#�������oN.��Xmw{�
��z��Ug�:�]���0�B�s���o3e��5oL��~Z!bh����9y7~�]�~�P��l�?A��.��:�������*v��l�'�g��k�7��;�C��֞�s�-:��Y����������� PK�j�f�  W  PK  ў,J               43.vec�e�SA���\�Cp��wwwwwwwwww	�)dX�Y���Τ�mD�����\�ȧ�)B�,�b�┠$�(M�R�=��H%*S��T��{j8kR��ԡ.��O�?Y4�R4ҍiBS�ќ���]k�6�-�hO:҉�tI9�5�覻Ӄ�������oʍ~>_=��b0C�0���a7R�b4c|{c���&�M����0�iLg3���s���y�gY�b��4E,���
V��լa-�Xo�!ˏ�z���V����L�b��n����c?8�!��;��q����9�ٔ�9�����e�p�k\�{��7�-ns����>x�~�#�=�Ox�3�󂗼��������G>�/|������?�C���PK?P@s  �  PK  ў,J               44.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��,�E]E�`v�u�m�L�����Nݿ���g����J׮�3��N
3�g`���:�Q��[�`�l֏.9�^,��H��w6֬���W�h�6_`��2Oe�3�0��dƂ)o�,f����t�䚲�s:7~y,��9�SrZ�H`�¢.<����9�*"�o�� �5m�KV&, ��G+9�H��/+��<�q�WJ4	MN]�F�(�3���pZx���jcV���=$ٓg&�&�����Ң �_���g8z!9r�r�5V+���s���P¸�b��&Ϥ	��ڧ���ӿ��H�w��|EݎEzO�.=]�ʬq�5��ov���[ƿ�-����� �5r_��_W�',)�����ԩ�L��ż`����?��G��r��^ԥ�ͥ���;���gǹ{���1�����\���������i/����Gl���W���ou�7�X�Պ�¦��2�		�7]]������f���gîD�L��.|r|��{Z��gM��ݤV�<+���\˔@W�&P(�u�#�{J�rB���)�V��2X3~]�;x�QV�B끴"�6��׿���'#�u�5o~��� PK(���  [  PK  ў,J               44.vec�e�Q��wN�؊�������������ݭ 
��Գ�ds���fGdY���K��0E(jS�Y����)CY�e9Q�Y��T�2U�J5�����&��M�R��4��Eì ��4�)�hNZ�ʮu���nK;�Ӂ�t�3]RNt�"�����'��M��/�F�7@d��P�1�)/Fڍң�X�1�	Ld��&�M�S��tf0�Y�fNʏ�v��|��E,f	KY�"�{�z%�X�ֲ��l�ۘ��&��-le���Nv�߱;ˋ=z/���r���;�c�8'8�)Ns���KY����/r��\�*׸������os����>xȣ�'��~�3�󂗼�5o<�[�w�=��'>�|��SA����E�PK���s  �  PK  ў,J               45.i��eT����`hB@�a@%�����.a��D�a@��P`@i���S�����_�{�s>��:�g���s��d�
0 �  ��<�^�pppq��pqq����(��	�@OI)h�h���x9�Y���韉r=�f������&���D�D4��4�,�,���z���a��01XO�10�1{ L�Ή����a<�������' ���Hx�����_5�_�E�M�" ��T�-.��`Hb>�em7P{�M��=����D������[""*&.�굼��LYGWO�������������������O��Q�I�)�i��Y�E�%�e�u��M�-�m?���!�~�O�&�S�3�+�k��[�;��'�g��W�7��� `b�O����q=���������4�ca��P�i�u{�*�G�21��,�}�t#�b^a?����߁����/���5 ���7<Lr p��$+��;Hլ�B���)h�Gx���m�?:,w��+g����w�wz�BF�>��R(��z���ka�����禄˵'�0K��	��8a�6�e���@[�fm�7x+�_��]8��(��i1��/�ݎ9G3.�nlC�hX7SbyVG�g���E��^?��1�$dwby�k>���b_�<�"�X}��*n|JJa�u��`���	�����,�=chƕ�+E���:��#����@ʷ�M&ճ嗢� ҅_q���zTLV7~����Jpxg"�+CY��[\~JZn�Lڏy5I6֗P�8�;��<��4^�;o�w��`Sa ą�)��y�|k[��}7��{�{�7���xAN�t%l!�s���+w{�M+���#�{"��+Ǚ��h}���t��9�b,7[/�$D��>Zk<�%+��*��j�{ԤX��3�̆q����i�_�|��b��?�~)t�E�^���.�Jn1�`m}�ec�z���lt�ޢ�$���p���?q`��+���
��E2i
�}o��}2Ɏ!��9����@o�����$f�N��]�vm��ӼDĒ 0,���I�Cn�r�@ĝrMYL���eVO�����`���g0�OW}��{h,ޟ�!֓�3ȿ����@���*Ը̅��8�8b�]tMb�#�w�)Ji�$/#��������E�G@�T�_�-C�e�W��@Q��j���,6�znT�IV!X�,���6Ia]��?�~x>ˬi�4�MoX�|����B�6C�8�UxY�uٓy��NT�LC�o{�nB&jn�I3:�t�T-�l!/���D�c�k�����Q)F_��.ע�}��M�%��u�~5�dk�d}nJ�mQ�V��Cˋa�ș2����cϠ�� �U��O�&���cW"Ө��E��6^pK%�%u|W^�/�!hk$�ߕ��N��p2�ٝ�F+$s�a�-�>�Zka}:�j���6��D�\f����7��$�gYk��^�'�h=I�A�/��*urS&q ��	c>����S0�5�VD�KM<��w�M�n(t�U|�W�[E�.�h%k�5�(��4����Nٞy��~&�Q����4Z��4N�].���Y���t�<�9d;DN��k�.4�	�w��d�b�V�`B ���g�7��R �=�Az'l���*D$��0yC�(���h��g��B�c��%~1E"��J��Ԏ�o^1
�����oS;��0�&�v�$i�Xg�&�	9-F'�?�Jq1�`Ɨ����t��"�+�d6]�RZ3�V�=P(p��\�W�	���'�P尽�q���b�=y嚫���Jd��+��;�tH$�����v��_��= h%�\���j�?���5kq�A�*-�~��kV��%�I0�|Ǚ%���׎?i��EÒ���I���@tk��N�8~������b4���T���>���U-�jx<z!s&"i��.�$�wWz��R���f"�CZ�vV�[�;�o���!���k�2V�P��9�G�n��&�D�ל��<�5��f��OrKw��6��m�'lm>		�5�������������Z#�֠���Rho��z�k���99�ޟ,캵7Ip�)k�D�A���O67��_7a�������x[4#��x��c�9���m��U$���*[%X�gE�y$��+ؚVi�/�SU�wɋ�U��K�����
N樔�\��Χ�ђ	��o]�����e#LŊE�h��a�!�Ng�����[ ���2BR���c/�K�A+h]����F\q!���m�"�鿡�^��Lv~�ɩ.���p�1�:�{j��!��.c9��`���C�%�iפǳ��q7�e��_3�t���z��PՋ���/J#S�n�}G6��w���"ȯcQ'�J)���]G=��/���Fo&�&��4ܫ�"
|��G�ŗ�Y�Wew�C�us��8�R������"�����.�\W�L�8�e��7I��zGF�t>G����q)��-mh|{��#7����3Z5��hT����D�o�˿����qxhQ�4�!�u�/�gdR~7��."������H�+:2]�&�e����ۓ�)�GQ�\Ҋ����j�Ƕ���z��liߟb74�
iL��	�x��ճ���Ϋf�3�%�(^�?�^w�-�e�(�!F�bǋӟʑl�Ǌ�	�O	���� xAƬ	�a�ew�L{Z��EM�;��<��g�/c&�� �դ0g������G�q�́�dS!���/�*�>8�Xl�~6*�����CRr�����_4k���_��,>:�Sw&�u���cv��,l���"b�:�)ovki�O3��7�P��k*���U�aiY���D2Ɵ�����%Z�]f�,.{Q���%q	i�o��Z�G���
�c(���MO� �j�>"OΥH�Q�Tʉ��; ��lr��Zv}n���s	𯊫eܖ���0���Qa;�Y`@b��Y�����/_G����,>x��bKF��^���٬l\��x?d&٫܌L�_������X����Dۆ'�1�0wz���<�?i':��C��̩ح�1���PS��}�C=�B�Dߏu=!��]�q��Ĥ<�X��ƷCfEu�9>f �
��^Ks�f�E��^]�^������vI�j_�Kp�ϻ �������M�b/���ЇF=�߷���Z�U�������n�
#V�	kڮ���t�q�nw{��֨����?�c�����{q�BӾ�]�pq��k"=���<KtV.�M>��K3Co�����������X��5�ə��/�x�/���ۣ�SC#,�M܍��/���8����R�҆��'������߶��8*Z7pH��<Y�g��)݄+o��'م�Vg���"�x�_��y^�/v7�$��-�l-�����$m���b���W Z���϶{�$���-���.�SK���M]�&1|��i�ϖQO�����z TXNh+�;6�k]����d�ś����W4���L��Kh� �|���	)���u��7$}/�6�Ƅ��
�<7&����*��V�k����WN5��}�p����xt}u�E�ۄ[1�BN�"e߮Lh��w�ͼ==!&4�t="�[���|-˖��A�襣v$��A�&0��i�LK�֫+5���rU�_�K��v�ܹ�wV����;�2���P����,v�$1�З��yhTY��y�.im� 6��S����t�'��"��\YsD`�aM�&ZBb]������p�(�EU��Y�~ۋ�nf'�#�A w�P)-1i��w^1�Y�w��̝CAZ�f�|�g���Cv�K���qg�mP%˻��U��h��6����!����0������F!n-u�ň,�f���1��
��_��R��qpO�ێ��y�����$�<��ȯe��`}$��Q~��R	��q�y����4+]<��W馐�=C�C�m�wn���:�����!%���HC�ES{Jr2H_SAZ�,�y~ǥK�B_H�'�1�Pz"��L�N��wo����]t� �HL+�R�J�3�;�r�����y]7��+fn�T)����e�6x���GA5�[���Q��.b~ʱ���ƣ������gZ���r�i>�4��79�Ќ�4��s��"������
���3�d@�N� YG��$��{�װYx�<~M��_'� ��$�и-��9����ӥ�#`� �N�YA-*����6������7
^�7�;���.�X��ze�6�'ݺ�7$���͗���qD=!�&D4���s=����`�m�,����g��.ZZ�,��Y���R�o�P�;
��q�ۺ�2��[��9�����Ad�[��_x�[�g�f�H��ذc1����Ɍ$���&��v}������3L_��G �f�Ӻp�hI��[a�c�\�Rmv�_��+�E����Iӷūƻܲo�D���ҥ���W��19��=�dR+WZ����3? CRz3��"N�|�gw�MGs��~�c��iNdv�EI%jiٻz��<X��P�|�u�!��2��,ۉ���j>�'����gO18��y��~t�pX�6�O��͑'g�Íy,q+��~�c��s�3<�0Lߢ�F����n�X̾�kpT��"��pU���3S��M����x�F]��H�;���	��Ri_DFj"��È��F�m�6��~t� �&̇	���}����<(�=V�1e.�;�ˣ���$��ߦE.�풖1`�8I�k�OFΊ��%��T����5�*`Y�qy�෷��ٱ��?H�Cj�M>#��c������Y����`U��r��2��؟����f���xT�n㟄Ksm
����8kכ�/�������sTm����=l�Z>y�[�*�9p"����'8�KB�Sc�Ӭ��S�H�O�,�W4�/j�j?�����dؾ�5Cq&���`�YR��U���r�y�-!�	E�a�b���A4=T����x;b%����b���\kk5��l=�W�4\_��Ŋ99f��ߤ����^�x�}���U� ������z ��z�ׂZ|f�[]�t}mB�]��-�Vh�
��HS~h����6�Z2�'O�k����0"-y`���Um��G���ZbI ���ݎg�I.���^
�g��V��li(E���U[��Yp�81�
�D��=�U���|��A�L�ӻ�P��pSJ{|Y��s<��d�h�..F�.�[� L��17 1���z�kR�n�Z}?vX UT����`���f?Ͳ��)/pA$1,�Ł���u�Ɣ��\�H��~�����*������y��{��P����s�������f1��r1ןd;�<�H7L9"K
��M3R�$ʪ�E�ߞ-BS]}c�*k��uD��BH�,����QO�$����ש
W���0��Tz3I�EW�h�?+������-�<�ޠ����{����&���4a[�t�D�7��N&�/şYP��jW�ҳ	��~��Oe�^��#��!�?Pբ"@� ��;O�;�o`4�&p&|4/9g��.�Q\���KUz(0�+o��?n�>�M(�c����d��4��ȃq{<϶��z'��b��)�8����S=����3�J`���J:Y���@�����!u�l�ӟ,��NS���N$�r3��$�%��O((�Y��l.#`�\V=}x�'��|�>F#K�]�:>�5�wjE�Gk���Պ�i���Lԡ#���_���%d"xb4�^�\�o��ʂ�u>6U�2�`Q��!����tF���E�v���]˗�-��&�l1;Wz*�)x�a��k$�?*~�6���z+o�Ŭ�R6�$��P�tx[�%�������$��f�� ����.�TV�Lª��GI��r�� �?k諷� ������ȭ>���E�N�{+1�%�I�� 5�尧�N�.����I8�:<�"����K.���$*�s��om�SM��b,S/}�W��h�����JqC5p���&��j���Y�'��z�֕G���[ZY�{��Li�M�B��:r����s�N���D9gI"bd,z��c���5A|�J��kE����f؜�ʼŌs��Z���jq��˹���-w��ϧ�H�ru�,?(lw�[�9[v�y��+I�l���R�cV�O]�2�:�DF\��$<*ij{h�����ȫ�Jl{�p�}m�z�i_�i��K�N�bђ�T7���>0<N�u1��{h��\��f���t���}�^�:�&g[���4ئ���I��ԏA q#8ُ6�n�M�WdIr/�?���Oх�U'�����g����S�wQ�UM#���Y�o�W?��s���P1.�H�^$�����<���ܣ!XU͝��[���J��3*�����B�8��O�����n�0��s������%Wӎ��lـ������N�bl���X�O�+��0:e�/p��U�WXD��N�-r5ɯ'�x��y{�����o�ޮJ��96��	�$�\,�^�!��ߛL��G�		r�iSHZ=�X��8��e�5�c���J��O6ը�*�8�')�/��.�	��u�xa�W�!�|�:��{�&|C[	�O�\=P0�����g���B�F�@�������o����K
�k#CnX�S%�5�Wv'œ/e�0]�{���L�Ī�6^R�p�����9���!�����������:�#֦Cbnp��*��Z=�uV��5�J
��w~�'4\�J?���"%\f���N7MY��C���*Eiy�ÒR�ڠ��k���k�r�.>�s�� ���m���F�F纤T@c#&�����*�b�s�'qTP���-��o�y��E%ok; ��~^)lo �� �/۴��p��V��.�s���X6�S��4ӽ��$��(��,Y��f�=wX�2+����T�lZ1AC��xL�y���9E�E�*�:��`3�;��w�+J��}n�WP��naZ�/ӊG�D�;�'q�iW��;Oi�& �1۟OF@1e�Ҥח����
���AE/ M�ߥoNg[$�?���c
���a��p�­��'�f���3�!ⴂ@������Kv��-H�)�����r���h�D<�O#0�����VЧF{{i��J�w�?uVE��[0�:�r���.J�v���i�8�|NB���Jje����|���b�я�r��;��s��4�~1'�'�Œ׷7���fb��� �`%6='��xP�a�fN�b	�V�W��b�8B�%�U����`<E���;)P>fw�܉¸��AB�� ��zq���z\�!� �>O���Z�@֡��ԑ*��収���_��U������i"S-��$��L+F�����5�)t������`�/YI-�t������;��L�E��ʾ�����2l�wsQ���2����L3}J�ꁵ� t�hF
�ܵ�:)�&N�����o�����ťT�e홳.NH�Y�'gF���Yz�d���C���+�b�D$[��ַ5�b�"ƥW���XI
�pҔG w��a���:�y�R�ɯ~_���R�حo��pm�9K��qa!2�Z�I����y:5���WV@�q.r�[�I������w�3�J5��f׾%�5�ahJwK��AQn�C�A�M*Z�H#�HM���F���+V����QU' tA�r[#�f��[Y�wCP&�җ�q�� 2��[�7���6��
� ��^���Īc?�U��P�Οurf���^@[��Q�.�k9j�1�Jg[7��%��ϐ�j���5
�KH��}��~l:!*���˫�y����n�v��,��O�����d����� ���ȇ�J�:����v'Lh���&���{���~���J���>���@��.��'A�^B*!��.���_^��{&�~���t$��u��쭅��y�f�rmtA��u�R�N۔��@(/.B׸�I_�D�T
|�M�O�p�zVҺX��}�i�.H׼w�'ʒeˉ�D���9=�i�K,�q�H��ܣcl��(�$p��;/�Y�����d9M�^@{�;KD��n��������1�C�h��D�����@�x���b��/�f�[rT��Y���w\/��uU7�NO����]��c�f��4¼G�N��0��}ȵ/��'E���������\�b�"'7՝�4�ށ�D�����R��%�@h�q�aJXm�<So�
���t-�I��̔�V�N������SZ9��#����>��t�����8�B.s}�FȪ��ǫ+��ݫhD��|��ty�	���@��<�����O��-��ט�K���-6��е�^�k{a'�Y_��G@͎��y��Bk���9��ˇ@"�GP�M5�[HmG�CEYy���vNx|@�]J7m/���m	�e���>�_iV(�c�"�+-phX\�ɡVZj,1m&�R�<j�du@����}��������wW�	��&0�o�)|�Q}�Afe*�v\J.�b�#��k	��v�vއ#8R�̅�b�*fc*������^�<4rd�Y�l�k�P�Sy��H*�+�9R���H-HpG�1���d[8�$�fp�J��r=9�OEM�SH>�Đ2���T%m�Û�h�-����(6z���56�H>�� �ɶu3�:-Hv3�l�}��/PK�#�"  #  PK  ў,J               46.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��,�E]E�`v��1���������?����l;�K����v�u_�p�,����8�z�h����N��}��湋����40���;�8�۰����g�z�)=��!5���l{f���j�,�y-��y��ķsd�ڶ��,w	��X��0�G.�]�q5ߗ:�\u�tqtW5O��`�vIӭ{�����)"P�bv���M�;ؿ,M37��X4�P�(�y5�w���?/�0f1�����L��*._"�l&q�g�z�����.n_m��N�Κ|bE����2���<�>������KL��/��l���`�e	�<���Oct�P�g%�cw��v�%���J�#���y��Y�st������/ۯ˜����`{��ջ>���=!���z�:�g����|5^/f���B~c���t�_/�[��g��9�K���4��ԙ����f?S:)Ӽ�M�����%z���U$Ё����B��K�o`V���h:��X�?Cu���]�.1����~a{������I�x�uU��Ů"!=���we�$۰дL����6s���+j�*�Ǯr-05:�3{~1c_Q��z�'�lA�=B��QLU��� PK���  g  PK  ў,J               46.vec�U��P���{��!������������w{� 
��H�r���ݦmD���+C�<r�(�(�d���$�(M�R��TH2Q�Y��T�*ըNj�I�r�ںu�G}АF4��D��0��f4�-iEk��־vI�u:҉�t�+��f�G�S��7}�K?�3��i6y��zC�pF0�Q�Ns1��X=��L`"�����7��t=���b6s��<�۷ ��B���,a)�X�
V�����լa-�X�6���fs[�V����d�ٓ���I^���9�Aq�#嘹����'9�i�p�s�炙��K\�
W��unp�7����w��=��<ⱹ'��<�9/x�+^�&�oͽ����G>�/|�[Z��+?"�����PK]��t  �  PK  ў,J               47.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��,�E]E�`vg͛�_���0��F��/��nfyo,��|�ݍ����iכy��gH���-�~%"������A#�#�?�YY��.��u���J��/�x�ħ?W_�z��4y�#���_�ꎽ���U$���ѣxxc���V���mg��T�Ƹ�̋6�<���F�Y�k�����Zw�D^Q��}���u�ъE],"���g�o35\�S3im����f�_�]��pb����Na���]����Ovq�j+|�K�����B��N���U�|}e?�����G>)�����{=R=p��xM��N=\z�[�߽څMҙ��̚�����e[ԓ7=͡���ڸ�'W+/b|�jC�s���_�N��*�*3^xp�m�J�װ)�/�_h�Lx7q���:�t=�mK��Th'۳0��Jkm��� PK�Mx  �  PK  ў,J               47.vec�SVQ��?T�k�m۶m۶m�d�v]�?���i�<�ߋ5��A1��W�,9�� �(����(�(N	JR�Ҕ��P�Y��T�"��L����_u]��Ԣ6u�K=����A��F4�	MiFsZ�ҾV1�ֺmiG{:БNtN���}��nt�=�Eo��7eC?s�� 2��a(���a���z��X�1�	LL�0��d=��Lc:3��,f�7��\=��,`!�X�����\X�W��U�fkY�����&6���lc;;ؙ~�]��n����c?8�!{�G�;��q����9�Y3���E.q�+\�]�=�}�[��w��}�{h�#��'<��y�K^y����跼�=��'>�%���{�����_!�PK*s    PK  ў,J               48.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��(�E,��`����ݖ�q�@�����V��:p'���7['~;Xt�p���$ۃ��i֛��}5�?�Ӯ�Il�_]s]E�a��NB�'_���C&�m��,i��OÃ����0ꉦ�N�9��������>�|���i����{�3���{���*�0�G.��3�$z>���G[C�W��]��f%�ʯ���ڮ첰i�.�=Κ:�&��/�_�k̹e�bQ�H�+�`���<��Xc�=���zJa�}ԛ�z�T���ah<�2/���������>:�U���p��Ħ�	��?�7RP��fo�vk�+-�}=ϐP��8�?Äy�*�.�Y�ڝZ���?w����>��}����)]��������ˀe�ͧ<��g�b:%{m'#�u��sJ��_��#t�.��:����[3��6eM���=땧�$�8�i$s=}�mW�1�:� w�TQZ�_�D���o PK� �ӈ  �  PK  ў,J               48.vec�ՎAК]����aqwwwwww���������I݇��LOGdY�rȥ y��)��FQ��)AIJQ�2����Y�
T���BU��,��ՐkR��ԡ.��O�?Y4�R4�ӄ�4�9-hI+�Z뵑�Ҏ�t�#��L��]���ܝ�$�^��}Sn���/` ���2��)/F荔G1�1�e���1Io�<��Lc:3��,f�7'��+�c>X�"����-�/��+X�*V����c}����(ob3[��6�����w���-�a/���r������Q��9�INq�3��9g����e�p�kv]w&7���6w��=��@�}���<qC���x�^��7��{#�����G>�/��kJ��}�.��'�"�PK9u�u    PK  ў,J               49.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��(�E,��`����L�u���ɤ�?������f�{����֎������Q��+ۖ?>�27����p3[d�
ρE]�	\��a%�4���J�W�&�f���BWW�k%=&NL�Zʟ���a�����&٪�V�u�N_�ԥ�`�\̩x�#���i�tBd��7\l��������ڴ�^St�N�����Mp���p�Y��H�����2����֊:���yg�L��V2�4�����'-K��ʩ���Q��̆�������3��𽎶�~L}�i��A��?O~_�������_�eo�������Ð��c��ɪ���I��֋'�-jZ�+͢��;e�����mU�
���|���D##�{����Yf����{����R�����Y��Vi,Z�a�B�>dw�o�g���IKaϓ��g��~~���z���jKw���Y䬶V�9��D�e���� PK����  �  PK  ў,J               49.vec�ՎAFѿg 8wwwwwwwwww�����K��X�d��ŗJw�DdY���K�(H!
S$ˍ��b�%)Ei�P�=��@E*Q�*T�Z~ճ���kR��ԡ.��O��Y�F�1MhJ3�ӂ��JY��k��Ҏ�t�#��L��]=_7ݝ����C_�����2��a(�Έ�#�F�ьa,��&2)EL����2���`&������"���,`!�X����}�ݷB�d�Y�Zֱ�)?6fy�Iof[��vv��]�O�ۣ����� �8�����1}����9�Y�ٜw^�"����r���w��oq�;���y���7��~�S�������������G>�/|��R���/?�O~�;�?PK�T�Os    PK  ў,J               50.i��eT������A	�i�s蔐A@�n��;$�Ia@:�kfx���Ɨ������{������z����&�XMIU	��
 ��[��5�< �� �������%=�KZZFV^vFfnZZ1Nn~aaav	)qAI^!a��l�������OE@@%�D�$����~ 	6�[@>
3 ���y���(�-��
*:&6.޿�b *
*::��hп8 ���I@�L��ك\0,� �E�a�Bw�/���g8�J*ꗯ��98��"�b�����UT�����0�����wpyy��~�����5*�[LRrJjZzFfVaQqIiYyEecSsKk[{G�����������ť�_�[�;�{��G��W�7�w����B���O��H�q�����c����H�1�0Ieu�,=Șð��pX�t�RXy��`�zu���&����"�_`��k����xh$ �^��$�|a�/����x�߉;�'���0Xm*a�e��.�KbƸ����t;�̬Z���&�Y�Fa�y�;q��w�Xᜀ��]�.m�P!��46��e��gOO2C�l��q*�G���=�{6'�Q�w�#�H�� "����ŕ��v��8�!b��d���>���S�c�(V�k�z'�NHT��x�T��Y�����wÆa���:	F��\T]*�gq=l֖�o%�Jݸ��2؁!����;��8�D���|ٿQ�V��oc�:�N��:�oZ��2�M����T>$����M��*�W�
�F@e۵�`q0"�Q���߄ �P�>���t>�x,�*r~>W�
�re��"��_b\9�Xê�s��J��w�'g	��̎(���I�;�����*m.��V��Ƭ!	�0|%�[E�P��$�=1.�C�0fW�ꗏ{���ت(�(F?,�	@9����Ա��9�Q	�vꯌ�D����IZ���3��ٗ���[�t⛮�����j=`��\=v0N��-�W��K�)���T�a�2 �d ��ҷ���ėh�G��k&|nbۂ�!\-s�~�'��Y�L����2u�N��>خ&���=B���[@+�]cY�܃B;�u��������Ujf2r��>*�̖ކ�"(s&�Ny��j��Ï����h\<�'����*n�*6���xsS��6S,��ֹ��$��f1!����`\���΋�=m����qP�wC|��_&?[���O�;(�	�-�b�?6ﾬ?���]8�g�j�5�D4��H����_ 81P��23�SP��3hCˊM�Zd�(��EkI?�_���.��9����<��Ή�a�`��S���w�W�+�N�!����X����6�����g�B���B)?%��h���.�M���[���H�b�l;�[%L�~l͈@�"�㷨��^�����>I^�J����Q����{������^a�>ʪ�`��C!hN�{�(�b!u�YT�Zfo���Q���G�Y��q��u�U�i,h}��(�Z�F�^y)��1�6%ɢ�-2S��ΰ����;o�ƫ%W�IA'W�>G_��2�����Yh�eރ6��]h5t!v�|#���Ǘ�)��~U�9Z��5q����'��ʘ'�}�{�I��Q�;��m��]c�]��\�t^~[���0��y�ϐv>�R���{Pt��oK�%��6J�EH:jG��p����Ʃ����`�?�i��v6��3�/9I{�)�1�1��,��Q�E���	z'J*b'9 ]`;qF�T��9���8G���X���梙s�E�1?�o�ώo��]���&bg�'��b���^��A֌���.�"X{UA1�6����5+i�o�9u�H@lC>n���,Jx����+x�~����Ѡ�r�.��.�ΐ_q�&��<�Z�f���uS^� �	��g9b��^DA���
Ij��B�ZP �n!W�cڄj��A�t�����l�vrV����Ts�����MWbN��>A��iO���@�<��3�}mԐ ����<]�mўTf�ۗ檕M���$� ���<-��3�������W�&70i��0=� }\�)���J%#�>�	��o��?�
��J��+u<>���,��,ʇ��P��ٶ|B�[�8~U�\% 0��!�+����=#�S�i;��*y^z0�<��'���F[`;�J��l!ŷ�GF-��[���0�
iǋd�t�V��RYH��C솀dў	�Dו���M�)���3Wg��sc3=\�1s�ʳ+�ؕ��{�:a?�G�U���q�4��L��ai�M�c2��
��:��y[��3=D���\����oۦ�7#*׬�����c��&��]oVw������o�׋I]ɓ>h�~�7fv��s�Bҁ��z`/	�*UR9P���U����([ǫ�Fte����=��F��~�k���>N�*�DY�>�=X��{�G���Jdl��mm[�v�qd�K���$>�K�|�Xٯ\	=^��λg �H#,d!K��d����,O�+O=�	�o�#
��咏g&��I�|���^:���l�.W8�A����j!^�Oݪ�C�6���jH�+�X�k7�����u���Ǖ��3�)|B�P;�n��X��FD�VJ���"|[�]��ǖ�Lt�D�]"w�(k=�J+���3�1��D��B�.���ީ`����3z�����)�=b�V�0@�q�Q)X�1y��<��;��7Q��C���\c�+�.�7�S��<����S�D���ۭ<=ќS�Ҟ�6i���P�"ژ#�����֖��@?	��ik���Ѥٷ��D���?�6��ղe���7���BY���W��I�D}�Ȕ��=�O�Y���?N�Ѳ^�M1j����-�AR��"��
EF���dn���*ߘX��j��D�N�v �%%��m�$����qM�'1����G�׻-�T֡�B�d�F"���e�� G��ɽ*�j[sh�gQ��	X�+G�.ùC�yH�V1w��|[?�E���^��l���d{[��MvE��&��l��/X~����l��s�� �o���&��o�8�S3��\��t�r(�π���rS������:�%L�G��˭���)���D�J���D����A�N�|�1�U�1HoEe��5.�St�K2�g��҇��P�?����<.R�o��f�c�Ғ�[�v��2�J���OoK�4(��X��-6V8����X�U$�c!13eׇ"�l�$�2���"E����vu@vߗ���z�\��G	-� nc��!�6�U� �S���n΍��ݫˡSr�I��Z�*��	��/_R'p8	�Ҙ~Kk��;"�1D��*�
e�<�-,	��n���e�@ϯ5�Jk�H���8ۅ���u���J���d��ɤ`K$F� *xN��NvgъU��7��h	XvR2,�$�U#%�C.7��jeCgC���H��IJ�Ek���iM��0a1"<|������ҟZY���7��G_�h��iG06��<R��Z�RZN��;5%��E�����4��o�M{����n�yRCn_�d�
�.�C�c�Ñ�/��i�k��YM����;��|���M�69�j�0�x��)��<p���$���r8Yn��,���J�h���]��-�^K���[���^�2�f4x֓֞��1�v����� \�6Dm����΍�ǽ������8���	��aQ=.

�{�uTy1'e�OD���:3{�a�d�ph�:��451���Kc��6�[!:�;�g�}s6�ƈ��ߜ�K�K����UU���C�ˀ� �2ZRJˤX�^CJM���=c�`+%�Ӈm�?P_@Z��KO�d#��hď��C0� 5S��|���+���C*�N�5l@?N�,�7U󿥞b"}jQeJ��`�߮0�_�"��ޫŻ��ZZ�^݊y �w� ��[��ڷֺ��� �D��ԧb��[d* 3�҈��&,?A����qVWQe���a�q��~qSe�Z����!�Y֕Z��U{�JC���H�3�@���u�/a����X?ք� ۆJ'9�w2j�3r�V�U�����h�XQ�~	Ǣ��ٛ�q�by3\�ѹ�d��I�����G����̍��}f��P���*�P�x�:9�`���hD�%��&����"�����*���屧
�w:D<�hp-M��)A�5��QZR%�3�7��R�W�-��-��P#���l�LAm��K)�)����9DG�S�V�:� ��A_�}�V,f�����%t����6��n�L"9un�8/P42��'�/%�2��F�T;���3�+_ �o�\�kD?g��ݬ�;OV�_]��K�����
��	���+��3���x_q��O�l�>�C�ӉΒ��)tEa��*W�i�,�A���R�}���[`��L�&!���E���͛��zOw��;��K��~�*�
�Ò��0�}:lT�s�nT��~�2'�""�lYE�����ba��a�1�F��2`�o1��,�Ǫ}�l��wow��SP��>�,�VM�X���ꄙ�T�_dϋ��+�h������_)]cM&cq��~��g|fI���d>�g`��p=#��u��,��F�
1af��K����j�!����*����������1�H��J����y�컪�ay�㯍��N?��Y#���ŝ8���Y���=�yN$R��!i��e�7peaz�8,U�X��H
S|GymҼm������K˥�������9��7�
6��y�
��d��|>�#}0������g���	/Q򠤺���ް�!�@���
b7���K��U�ڏ��t����O�~r*��џ*����o�#�(h����"7 ܈����Rv,W[�h�@&i.r<fnj_x�h��>օM�YS���%�ʡ`�*�t�[�y!��еW_�1]�U��c8�v|0��m��B����g���t�]LW,k./�\S����}NV�̚�.�Lo��̈G37�bm.��@N�2;���z����LY��Ԛ;Ҡg�&ч�p|h���³���D�:�^�*dM�E�F�8���J��u*\�tBv�^`X>��l�r�
_���C��������>IL� }S�~�����WD�Wb%�B�ܿ�)�~'6NBԈ~��G�gl�ofWAc!8�_M�߀���z0��'�ګ��V���2^_�G����p�٥�6��VV7�;Y�|��õL3�Lj���`K��\#��&���u��s�<]��{6�师x��j>�<�<"&�a択�m����r�Ư�L��������r�z�iK�o������^|���}��Sy-/��'6`�B������lE�Q���^�F5d�O��Orxns�̓'���!U�u���^�$y���*��!Y˴�,���cC2�rA�St׻R�%)���4XA�0V"�p.[�&�\�T�"�X���Aw��CLZN��ׯ����]�?�m�
�E���A�P)'{9�ď���ɭ+`o-��Ӫ��8c�۱�9[?"S�f�?��]��
$����4�~��ǳ��0?�|�]U�eu�	㟝ޱ|����[E�͸�����- /�֥��Ð��'.L3߶��kI�&��Ό��C���� ��5������ȕ���`�\���W�D��h54�;�'��s�m(&��Ӯ�(<��}��r�'�v*�SM�=��=B\��
�� �`Qщ�<�0���ٓ��/�_�¸P��z��*X�Mby	�S��k�^��}���@�Z<�e�#�{����pY40�U�C�1�����!䦒�g%�OX���}R����+]�)N�4/�u���~P嬐�h�lm�i�'���c�[:�Q�y$*�!L�����M��	o?�4p!�~�i�I^�FA�����+"1$N,	�u�A��.�	(�*,����N+�	*� Ow�]P¯���ܱb	ٴ,*�����54�X�M�.{)�j�0@e{�D�IWp$ر��ur��ϊ�����L�Y�����M�\���)�M��g�(�?�c��][�ͨkxփno+g���=5�[�<Y8��G��e�Dj��`���{�Js^�/6�Ű�b˾�?��$N=��%UE_e�QQ�;��tyѳ��Gb�X쟃�ض�f�"�4Tl}l��2�޸�il�Pn�Y@���j�ɔ
7`�a-p�ΉOgv��,*B��9;���Ƥ��~����X]������?|�bd��yQD։�\x�)��
C��5�)�t�E� '����@âR��l.}/IIg'V0I����G�T���v������Ѷ/��O�8�#��ӯ/5�9�҆��]Q:����:��n:�-}Ma:�������{p����4�]�e�`?�7�v���PB?�k?����|w�2X_u�H���{� �8}�#1^���Q5���|��:�)rv:��ɸ��K���ҽ����7�\j�o��N�r[��5=�\��0'��f��|����:|ǉ�P�a&�[�z/VB���%��x�O�/�����(�h���U���������݀2?��9��s���7�u�TF�$Ȱ<.Hӧ�FgL���ع�<I|D������E�	��݌Y��ԝ�i��xW}@���㕈$��v�m��3t23I�H�����P��cKTh��P��I	گ����'u�z�*��� �*�����E�I����:��wi�"r\2�z���x	�=��m���%�:)��� L���E6�W�c�noQL�!%v��ы�o#';�8��,��Ȳ�2PF�1F^�{!�+��_u̘ř6�)����ioD��Tă
�iۄ�Ft���Ў��yL+.�ǧK�+#~��aaJ�a:4Ɵ��y1oJ���f\�N��֡�5�π���!�y���,u_�c�Ug�Jr>�b�
�����~���8"d��B����\��μ���X��*b�)�e�����p�^E��P��2����n	u�2W�#��>l��A���>�����D�!�2/7�I1�z�M��?�`4\����e9쭵*�+T�d��G��ex�5&˼��p�X��1ن��X���Ę2%�����V*'r�PA�J~�jG'k�|�~M�K��H����򚴯U���}C�J�����(�\X#�{7bi1�ɕ�x�G}���̱�(����Bf�E� >0�ԗ�$�3h����S��  ���G˖<f�H�P�d���7��g �2�C�zpj���d��E�>�aʰ,��gv��ȶic�M�v�b��3a��b00�0�j�]/��EHT�/(x
��7c��L�-y�ƕ�+I�U�G���*h�c����2���Xz�Y%�V�?�e��E� �Dn6�'{�̺����4��pP��(D�^�έ���=�t>9�aK�,ϔ��ȯdd6�(bD� I��\�{IҰ�����V�3rv��o��9�&�e�n����ʳg�s��H�02�q�A#]\�-�J��'���i��;��*l���5�Kk�MT��H�]�ݿL�Q����\��>:`�ȑq�����n�2���Mu�"f:Y�$4����>e>G'����:��q���^,���S���*�GJh�%��,�I�'���b�)}T�C.9�ޖ��l�G��Mo�+gL0��
"!;�=>z#6߲4H].{W�׵�7"9j�z�ƈ��cƁ!/q�J��ԉ���C�:�o�%7*A��j\o	�~�I�b7�j0�@5���/�������B Xb�ƻVAI�0���l���ԡөh�&��z��[��A��L;f�1�<����\rb�6�?G�We��wA��:�8q.�;�3'Y͔�(p���#�D�Ԓ�{��T'��t���8v�hmi��	�+�c�������J�-9Z=�F��V]T���Z��-n%���2y���хRM���dH��Q�S��8Y��'�m��T�.�L�4�����l�.��vy��8�a�F��^��o�QZ{��^A+�:�cE�s� �L�z�h�������0�p=?���,������]�2���W�z��oJ{�J��C���
�-W�����;Q5H9*�;�Mq٪��_(����=�#�d�'ÊU��O$����K'O�:-���+�C�΍+ɉ��`��\�*�~���@T�eL��i|9�mU���ֹ�g0��r+8�c�NS)F'���A+%�!i�$jI@	x4�Pnz����3�cZ�K��֍T!{��D�_�P
v�B��<	����r��W+�/]c�ip����}��/{x�~�E�����U�Fר�������	X��BR�2���n)/���������x�ev�-p�3��*��(�����e�F[��n�Z`jfQ�HX��p��֔�Ԩ7�^&���[�L�f�S�ϔ�Tu�i��%S��>uWS��[AV���J/�QÏ�+�c� ��x"�a�.��ɥ�[-�R��������4�^�_ח��L����"΃���b �h�=��o��71����([4���|���g���5���N��k}z/��&2����#���%���D
�_O�����K��d�J	�"��w����\�V��2��oX��_���r+%Ͽ�PK�%#�"  *#  PK  ў,J               51.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��(�E,��`����^%�]���(�^j�c���[���ϰ��K��l�7���p�~����у'4��gp\�6S!MV$0�!�U�f�8���Wfa�A(���v�";�v���~�I��i"[��ݽ�B����c��¸�^,�J	te�#{��]�T��x}m��3����]{=33����{�u��mg9Z�[��������\κ��-����&zQ���@�:7�Z��=�̬�1�V��zb�A���ئZ��U�PhﱇM7c��^[ ��:�n磕FJ�\��l��K�^�N}|�MLk��W���/�7�u=u��WS#���d�5r6�?�����L�#የ/�[Z/쐙�DA~��S��o�6���.�+,����;Rc��k/<���r����ꧻ���TI�]�"6u�tѶ�x�;�*RK�]�������W#󶜌���q����N[��,���z�6��X�w�3�n��s�����DZ.��ʳ����޷�ݷs�;7��P�g��p��W�k[�)��	 PKG�M��  +  PK  ў,J               51.vec�S�Q��oڦnS۶m۶m�v��6S���S���j&+��x�'�LD���'�\�ȧ�)B�,7�9�S����4e(K9��wV�"��L�R��Y԰��kQ�:ԥ�i@C�FY�ƺ	MiFsZВV�N9�Ʈ�nG{:БNt�]Snt���=�Eo�З~�Oy1�n��`�0�ag#�Fٍ�c�8�3��Lbr��b7UOc:3��,f3��E��X�"���,c��Vd��R�b5kX�:ֳ���ol�۬���mlg;����'�������r���h���q}����4g8�9��\p^����U�q�� n��ҷ��]�q�<�oxl�D?��y�K^�7������G>�/|��R�����'���PK[&��m     PK  ў,J               52.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��(�E]E�`��GL�rn�����ck+v�9������o�6���|���ymn^`�hwߋ��uS�=ygl	t�RXԥ��3�y�뻅N���ɲ\9�a����������Iӝ`�{m���a����j�}��hFS���Q<b1{���y��1<��]]o��j��E���q|{ ig��mo?7��XfV��޳R�& ���g�U;;l�C׌�}��1�3=&پXꋿ葵+�j��)��V�"W�o�'������2��_t���XԀ��O���c��ҜyE��v�d?S��VV��ëNtq3\��x�B���}S�&���~��וG�1�)�V|�b��.�g��C�o�������$�=��%�q���Zs�F)A��
ܿ����y�{��*����y?�g	�^�m�g�v[WW�M-�y+�\�����������=��X�d��㈣�ҋJ�-��;4��D���l���t��7�q��󏺒�/�3쵎�ē����)�M�ځ $�ʀ��]�[vZ��۝�m����_�4'�r��0���|���B��޹�Uq�/{������Lw�� PK�ғ�  \  PK  ў,J               52.vec�U��PЯwf�����.������n��]��@�?��H����N{N҈$��O��(BQ�Q<�D	Y�R��e)Gy*xOEY��T�*ըNj擨eW[�C]�Q�4���$i4՛9Ysق���5mh�D�$��ށ�t�3]�J7�����=�^�������fc�� }0C�0�3���Js1�n�>�q�g��d��M���Og3��l�0�y�7�=�Y�b���e,gE�2��*}5kX�:ֳ��lJ���$[��lc;;��.v��no��}�~p�C�G9�&q��~�S��g9�y.�\�����r����f��[v��;���y�C�8�O���x�^�׼�;�����G>�/|�[�����C���#�PK�;�s  �  PK  ў,J               53.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��(�E]E�`�-۝=������?�ژ��?7�2�o���-�`�YD��4��ܬ�OI�����^�ܵI҆/u]p$d��o�b�9{*�d���V��<�v�_΃��u�<���W穾b=�ʿ�5��@3��45�⑋�E��|�YTҺS���B�H��=C L5v�;O~%�m={�'v�����!S�\[6U$0�`Q�1sЋ��{p����+��襥�Y�o;�*������6�(%�r9��5��{�L�1���V8��Kr\����ϠitTP��R�B��'��'q�?/��)���˕U$������b%5.��~���/cJ?�;�;64�=|j��F�sqaLL{I�������wf^cK*R�5�e8�/���cK{ʏ�?��β����5�ӵk���H�.x���z��o�|�����y
:|���E����ע��kK�_)_k}R4�Һ����l���pv�ז@W�du{�0v}~������y� _M��w�Z������[�m���������sYՔ�&.�pU�X�ŀ�_�z[,�rK5~j�q��?��n4�Ǻ�m%WeyO[�%���3/{2��G-�m���� PK��a  f  PK  ў,J               53.vec�U�AК�����������������%8�S�i���}��t�'"����G>�(BQ�Q<ˏfIJQ�2���`OE���BU�Q��,̢VQ[�C]�Q�4����d)���hNZҊִ�mʋv���;БNt�]�F��=���܋���/��� ���7X�P�1��d�S.�荕�1�	Ld���T�iz���d���\�1?e��=ʋX�����`e�X��jykY�z6��MlNb�7�*oc;;��.v���z��\�p�C�G9�q�;�wR>�i�p�s�����y�+\�׹�Mn�¸m��.�����<I��3�9/x�+^󆷼�=��'>�|���K?̟��w�PK���n  �  PK  ў,J               54.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��(�E]E�`����z�%�p��{�9�Oп����g�tM%�MW��)'~5w]����Í��v��i[Gy�Xԥ��*�K�N�ε��Ϫ��U�]���R}��<}�sɿ�!Qw6��W�Do|�)��V$�g¢.�Q<b1����/�VZ|�9��ڛQg{;}���<a�Y�e��	q�_��V��>�*T�D�=دKc�D��1���]O�ʧ��� �Ztl���3eJS����b�ϰj��D��E���v�:�!�Ͼ��Wޝ<��u^����I\_\1�g{R��φC���~�����υ������̣w�tO	tUlœ���~eI���g��9��x��w����ձN��l�i���ET���g�c'<'<���O�qU�e�������ÿ���ߪ��t������=�/�g�M�k�;1��ʶ��X���|�]�oCo��|�v��<^m��oI���&v��PN�om/�2/���rz�;�?�7V�?m�q�-g0jt4u1`�/K+�FNuj+`����]-M��z����b+>.�(����g�Z�e_��Em֍���o PK�}���  A  PK  ў,J               54.vec�e�Q��g�9�������������݊����?��]2,���f3�e���#�r�0E(��E1gqJP�R��e)���
T���BU�Q�o5������C]�Q�4�k��h��Дf4�-iE�m��V��=�H':Ӆ�)?�y��=�Eo�З~�O1�n��`�0�ag#�Fٍ�c�8�3��Lbr����zә�Lf1�9�M�|�|���,b1KX�2�ۭ�r�R�b5kX�:ֳ���wl�
b���V����d����o���~p�C�GS������9�Y�q޷^p^����U�q���[�6w��=��<J����g<�/y�k��w����g�D��)�7��w������PK�n��n  �  PK  ў,J               55.i��eT���J��nPZ��!����.Aa���GzHA��:����{����n|������:�������<�=���+�)00 �� P���qq��@ >>�"BB"2r
Z&FZzzfv�̬�l����\��"""L/$AB2��"B�9������j!z��g=vH�0� ?�0X��X��} �����o��00��qp�x���6�?`b`aabc��`c�����Iq�X�qɵ�Y�)�����j�)u&�م�<B�	�QQ��r<���-"*&.!)��JIYEUM]WO�������������������'?�Я���#"���SRӾ�gd���J�~���7465�������CS�3���s���7P�[�;�{'�g��W�7��pa �0����\���0������������RlA\2ym�{wrV�`<
�ļ�n|6a�cJ+�I�g�"k'�A�o��;���/������DX���"�g�7O�/�ˬ�ML����]�X?��m����>v<���bssR������,�_�}�Ad�}����eF`)A %P�;�/�v[�]�Z�Iq6�Åy?�9�S�tv�X-��L-��uW���I��:�[Oы�W���x�䎠m�?�s�FL����5�o뵀W���N��g������c:�
�:�g�P~�p���s�PP��2�,��OB�,\A^z�paZ܁M���s�������7�Ģ�=�����q$g�;е��i���6GP� x�4�zV�J����Q��5	|�X��\��U�����<(�t$�x_�;���*nGi��ɉ�C���*df�"������w�9/�@��y��fq�"�ߡXa�Nz�d�gz���%�����*�0��E�>��J8:�8��T�f�\)��d���p m��u�^��i6'ZgQk����7
��/<���˚ߕb�{�ʈ��'7[Ųq{[���������c��F��j��X��Ҙ>�3�!�|��f�]�)g�*��#exc�x���~��K;�g�!�U~�OL� �#c=�<�xm
��y����t�x�P^�=����Yx��[<I=�h���2PgE2<��GWJ�o�(&!&tX�R��.7+�!3�z�P����z������	�S�h���|� �d�j�����D�LUI����ĕ���㵿a��z����t�ӧJL�:y;�s�է��)5BF/���6�7(TG�����6/
���1`̳kͱ/t8�!��|�$�T�F� (9�{�t/��W�K(n��=q�z�_7 �K�:�b��L�t��Kf1H��0�"�We�X�{�Pw��5��k�sM���Y��o<�������ϴh	6C�q�|ܓiX`yv��x�"&�����?d~h:���5�:���4�����o�D1�G��I2<���	>mq��cν?-,L���@^ljk���я@!��M��<��kQ ���ڹm�ĺ�Y&�+�<-.�����0�P��݁c9�FW3-�6�`�z�V�D�K5��Sm�1��Z������+*���\��o�7}i_�@;3c�������$�KV���� )�YL?���f���M0�\�rz����m].�qA�W�g�xs�-m��0�7��D�A{������FP@���KABs��<���)���n
<��}�̟�w}�=�Jo�`�=�p�p��l�w!�����>��ԅ�W�7��8����k	�0�r7(�|0�r�]z#}�x�����⨵y=�3�*�MF�\''��^�X��T�:��3)�\��ͩ U��&֗��!�. A�yټ����2�H��Q�j���R�|Q���J�8���6�&h�A�!���0p� �N�*S�� ���A�y����YahO��=˻k�7+�)ra�����$���J^�w�����:�o�6��N����jg������]��E��R���ܝʾ�t�n^?�m��48Ǭ:�oَ�ZD3�-�9�C*���Ҩ���v5�x����v��D�'/��XT~��#�пI}]b	�
r�('�M�B+�ðH+�5'��|dG��Ҿ2������{%�Z!����Eaf^y�G �.�W���6��.t���hM���h�>�Lܤ$��/{Q|.��?���{jt����,b�ǰV�I����MM���W��eG犬�N�R�%�$�h͍������Lw�%-<�lT�g�'��.e���l�i�[F���}�K�Nʨ��2�/���<NŸ���sS���~��^�k�s,�}��<���)������{��S1�wAx���sԊ{�Y����W�L�����{��6~� b�M��P]4�b#��*-g�κ�~�<�E�oP�:s&[�H͗���Է�YW1lB��U�@��,qj��q�wG�U��\�mP�������L�m%Iu��v�vi�9�F��q��^l����Y�=��Sn�<$y�i�K�̺�&i��$k����|ki{�sU��r6Ƀ���D�A�z��]Rf���H�e���R����*��jR���8ˌv/I�a0��2&Ih�̖1 TY� QY��ᐡBNj&�8!u�T&�@$���0�^�=�$�� {>*;<6��&�&��|���5z�Ɇ�+m��"��2�9!�O���
WeM�.�}�5߈R�DPˤ�@fZâ5�Q8_�=*���Y���8nS������	�B����sJ�y|�G��\p��*��KvY?xQ�����⏂@�\B���=�u���c�0.d���P]����Y�b�GJ���?����4���H�f�5K$�f5�����}��Lә;/�gr0��7���o�����b}�	��3��R7V�_�kͤ5r����0��߁	4�
���fЇq�*6��ZRZ��l��hx��TW�B��\��h�`��:!-:�^�F6�T_��/9Y{˂Q�W�>g6�~�ϲ{tT�p~���Ɛ@64jg+�FF�75�-��o�&ʫdZ�&*��.�f�0�Xq�>�]����N	�u���	๛[���΋y������"���4@]}���)�V��ö:i��{�MC�P7���%�q��!�����%�<�}5�꽯��\l[m�lޡ�*���oF� /�Q�[����(�Xi�왟��6�[<��!5V|X:^��Ɨ�� �}c��� ��X��J'^Y�%"��Q�=�?"��';4��� 6���&��3�
&�,K��wG�����en4�Ӯ�[��A�]�5�9���:E���=�
~���J�A>�]��ͨ����i`t/z���H����km�����.|]T��ɍI7jGt��!x���Q�����A��徉����#B�����[HM)�+���eS��v�I������X(�J2�I�s��Oy>u�:_&���y�0����J���hB.M&rcS.�!���sY^6�@w�.��i�&9]&�� ĥ�.E�nM0S�$���MLu�����Q�2���P-#��|�H��8�#؝�����1Iς��e�~:g�����IGq�G�E���+G\l�i�t�������f�����!J{U\�!�m�ğ���~�t)���̫q,�5}����J0��1x��<��xS����KOL1K�^G�@�*��|-r�ٌ������Nۺ�"��z;��r���R�M��������i�9&��?:��݋`��ޡ�HiyH��v�vMo±�����2�t	.P���4ࠋ
2ĸT�U:F��z�	�t��ӥ� ��>���P���31�fǞ��Vj�c*;�l��� ����%+a�Є���Vr?� ��2��Ǔ6�ΖI v��Ľ_��Zdh0�iBsN�*ڏS0����q��|�K��]��sF�~�����S�T+�̕��H��U4�[6�b�6���u�2�;*��.���6��쫶5������������A�r�H@7qԤ��9���Y}�~��+�S�,2���%��!���D��7ml�%F����2��.j.+z�`1�B��@e测����AP���%٫���y叵Ij�$?�+�[�,���0��5W�tCN�rv|�=�A 6�I��V'�A��VJ��߶k�ϐ���`�:^]�>y�$,����	�u����_k���܂��|a��d�ANu'��?y$���t�6�����B"��}Ρ��.�3,u<����ڍNs�iv�|�����T�`��;�vFx�pV����Y���^Zlt�f�g~
�ګ����|b4U��Ah\�i�D۸�v�K��R�j�	���J>�7GT���xz�KhHEK$�#��JSַu)گ��&��G����v�h��d�J��9ꬽ�%����ӈG@d@��1����������!N;��Mb���
�^�H��.�9�F mBd���x�u��ҹTSd�0 ��:� P-�����x� �I׃�R��&���Qv� ��(P�4�;=ӟk��(οlT����6(Bޔ�cy��n�Jv���t�
wb�f��5Bט��rNạ�2�?��.z�˖:K�r�����6=���)�uD�\�9@lfܳZ@�ԙȟ�_F/�;'��� ;j�rԓs7ѓS���8�6��UZR�e�m��=�ҧ�Pz!��܌J�Z<�	����x�VV�Ǻ���c{"j�����=g��\��	aw�p�w����Y�Y�a<����6��;Rsb���ٺ}��A@���6i/ɖ�3���A:V��tj��J�5��sR�"�?o��̞H�vn�kN/�u7Ĝ]`ks�P7ؠ?-�y=���С����>V��2�"�8dh�#���q<=E���=�M[RB���&Oj6�]\�>�U�ST^����&���I�6@�U]����I~:ϼIb6��(�� �Ҵ�m�[��{U{�j�exp��Wts�'B�
���NP�A��&���%[���~�}�0ER�׼C�(ҶG@����#@�i��'o����F��a�1�&ͅ��f���I6M�_�=>tf�qie��+D�����G YE4�I��A,�50it�׷���,>K�c���4Y�9eFo6����ۦx6X|�ޗ�䣰��<�K~��͍<l��>�<���C��K6�vf�ۆ� ���L�������R�b�='�W_ߔ)6k������ '{9����nLxu����{jhO��YƲ|'$� AuRR�~D��W(�E����jliJH�N��e�+cE�\	-\�Ⰸo��LW��|�-�HJ�+.�o��YP�B-Z��i��Vd<����DGѳ��^Y[�a�)��O� /��M�s�a5#/u���`�f�b��b3T��?���Y���iR��z�y�k&���Om�E�W��QF��ýPv�DenCv�����~�ѥ���k����97�G�G����z/�iغ�vf�1�y羛�UUڍ�lk�iK�g�ؤ�-�썸���M��3�?��{3�*
L����|���?��fF�|��W�$�Q��OE4��Ԭ��Zi�,���-.��ܚ��I��b�J'���C��!�7�7fѿ��)(9:l��(o*���x?��+��deH���W9de���ʸ��m�''�U~�-zü�_|�J�d[V6��7l�)%>�A�H	�&��n�֙
~�nK`Ās�0> q��F>�$��=��� mgL5�����8<ќ1$�k�ܼmA�mC����+.v����f�_����)ƀ�B�����aTcK�Y�����OBڽi�.��=0=.R��GD�oa�/�l�J"'3-�� �Yw�I�Ғ��P\�G�@��P�.r��&����غ�F�`��L��Ы�W�&D�~V7~��=oJ��Fh�v��ϓ�wO}<�^uY�M�ڥb��5����X��Pv��	�Zs"0�ّ�Y��D�J*��Mޠt���X��F��>6L���@��c;DR���6p�y�Hr����seW��՞lUS變�;�Ʋg�o%��9��7�U��'�F�P�E��I�>6g`�Z�!eƖֶ�V:����c��*�Y���u��7�/���K�^�#ղRY��\��}�I#�L�ٝ�F�:�蘼��V1X��:�ǽ&�S=�*9�Z;�{���uZU���l6�J��}���B�)5|�ͣLR�d��Ķ,�����Q�v�c��{әz����E��e�����By](甋;���O�~6��#���kk����6VU��$O��i��:CG�@��[.���w�}�O�	<`���Bib�\����CV�g0n��@�����*�����Q/Dɗh��ܪP������{�*߂F�����6���׳vSΛ>���\�J�#��x���d���Pau+�/ycR��y�qwO�����R}[�O��ʗת�aSx���4OmǨ�]VRm,�ϋ�:Eq׹�Z��Za1í3����uN*oi^�fh�d�6�\->kW��fk$'\(����)ٚ@�a�s$�Q����%f?06[���_|�z�;���)��R��n4v
��xv����V��١�>��<3	�e���(`;+��\�p�%<���S
�)�����VR�WՇLJFF]5�_��&b�����x&b�n���3#o!_���bVR��#|���{љ�}I�~�jJ���D�?���4�u��Cxc��̗�ɞ�$A�����bo�<�m�6�&�\Ū��d89�zwh.�TģgIY�k���D���o�/5���!��!�ZX��r3W�f���ʫ�N42�0�p@2&�L:��8;���4yp{�%
�ۊ��R��	Mu�I��ў[�"��Z��3Ç��O���F�6�!Q%e�������4x �u�sI��O���B�_�/�2�K���s���6�����8	�q����c�i�pZ*������	M�6�gn�p�Ґ���G��pk!M�RS� 6�&"D��A�0��j����<MD1-|�~�'���UL�V*�zUO���j/O�<��r�~���R���f�د��)��Rt@���;&$
��Y�,8�;��}�*>z@ �ճ�LP�h���}��&�S���S���jD�ҸK} ��9�����X���0| ��o�5NRF�AC��ͺ��/lDf�Պ�c����!�q;t���o{%-ݑ���o-�s��n���3k*�dbe\f#�]�n�D
S��&���C�ld0�?��YN���F/�
ܬ���򌟪f��1��&�V�꼹s2U��O'M7����כ�c9�?8�՗��B��:���eA�LE^$�s�*K[��*ꇟZ���)�o���z��<ܞ��Z���%JB7�T�.�#}u#�u���W+m7� V"���O�ln�R^���н侱J��>���%�kDW�A�LH�r�9�zc��731ts��e�w,}�����x��ٌ�"Έ�dI4K�)Q�<\9ʠ*UTc�m�I=����m,K����Z6����<D3�������0^;(��Wf�X�P��ޱ�V���ĉ�*��0UpKn+'�i8�-Ȱb�t̽v~��ڔ���j2���f6�(���n\�:�$�r��t��I��M?�˿N#3}Q�v`�0�B��>1* |��fO����|S��.ӡ��O�A�>@U}���+^M�2����F���;�w�bu5<	Oc�S�~xa=�Âd7_�>�n���sp|�w����_��t�(P�U޸�2P��J�*�g��d~Ó�a��D��
y�D���I�]�4�s0N�=�r~�-��9W�����H��vVa�*A��}���Ŝc���c�=�#�z���4>3<��������A@E�G��E�U�'��w��~	�7?�{�'�w��� ߣ�#Z���`���.��x(��9�&��~�(��{2�aS
d��6�h��qQ���
p�p޶��t��������D1��i�c�~����C�FO��D���K��`��pj��fnN�B�M������6�@�W�s[�
u��A�f��0YD���u�O�AK5�67n��Ousӥ��VZ��S�3�|I�ԏyC6���Y�J�6�o����n̖��� �B�n�����~�b�5<,&�71�8;t�[��~ؕ=[\z%d�u3�.lh�>}Yc9�W��Jv�u�E��v��x-3\�Ƃ��V�{�.E��Q�dL��c�Wx{�k�he��eb��p!C�b�d��VrR��JnƄ$	%��W�JR=;�	c�^�k����N�M�t^��!���у,��u�}�Djc�L������Oa]�g\�,a$�U��-�Y��IW��W�T��eR��f5�E��p0TY�	�>6�_e嫘mӅ�%Pj$S�����yK�鿏��= -y�̌	9�@>1�|�����@�v.�s��UN�z{�BH2��Q�e	q���IGZiy|���є�@�4�{����NF*m&~�[$F]��ܜ�	��<��e�$��*�����LE����Ԍυ�O's:Nv�K�β=0���u��D�d�PjR����p�$��1G���H_��l��8�`n��i���U\/c�俒5�*;�V-Y�|�g��!���7/���4�]��T���<�9jT+�>w����P���1���{�_���k����ֳfV��ɸ޼+{S\�������ʑ-�L#�a��~��Eo$�?���o�9�dt�2��%$ॾ���MR�y��=t��8az��_PK�gξ"  P#  PK  ў,J               56.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=��(�E]E�`֎u�"���~�r��Y�>J�ܟ�P<���MG�B�e�WJ�{i����H;D]�������O��]E��45��:���+|b��(�}A�k�Ts"cPY���z�9���!�I
)�L2B�/����2��QLo��7���E,��Ȫ���Sr�vk�.�Y������A[{��O$��.RN_�c�­��;�;��w+�Tǰt�>� q8|QE��ԇd�5)�^dP�3=xj��3<�}vS\'M��L�<��p��W����`��xs�m�ocj?ϩ�^UeG���E!e���sR��g�?��]~���QL��'֖���K��n��s�ߦEL0o�ߚy�����)1�������;9�޴��PqTU���9o��l<���뿖�����i��lg0�ύ�9��(���	����s�i��&+�EK6,��`����C�u��.�z ��d)��'{±����G'�ݨ�.��'2}�v\�7Y�;ѽ��M PK���    PK  ў,J               56.vec�S�Q��oڦnS۶m۶m۶m�M�^��9�]�de��7;3��Ȳ��K��0E(��D1�┠$�(M�R�9��+P�JT�
U�F��,jd���Em�P�zԧ�e)�&4��iAKZ�:�D�,��nG{:БNt�]Snt�|�uzҋ���/���b��@=��a(��F:o��h=���c<��$&���b7UOc:3��,f3��)b������E,f	KY�r�Y~�ԫX�ֲ��l`c���6�-le���Nv��n��^���� �8���,���'8�)Ns�����q��^ԗ���r����f*�[λ��p�{��y�c����~�s^�W��oy�{>�O|�_#ŷ�����/~G�PK��3o     PK  ў,J               57.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G/�E,��`���2�&4��Rz�0���|<��9���b���3�\��D�=��B�ݜ�/+���H�v	mtaţx�bƍV����0(~}�G���u�>�M�;�����_�Xg��Y~� ��q:��a;&:O�:�p��SǓ^7L���.�B�͖cb�k�'ϙ���g�:����l�w���ޙ�e��H����H #���V�&��^�܆O&�=�r���grj�7\M�)5�3����;!�s��g�?��;������u�m���J��;���ʸW��/�8��l���?[�ue��l��ȵ�~U�*aK_DꙜ��.܅���������6�iN�/�����0�g��Tf�B`�I���g�-��H�)+�!�ʀ�Hm��\���Y�-�����<i�f��Z����R�+����ޢ�Ɂ��ճ��e���	 PK�� �p  �  PK  ў,J               57.vec�S�Q��w��n�ڶm۶m۶m�vR���S���|������L&"ˉ���.��#?(H!�®E(J1�S����tʢL�EY]��T�"��L��ɢZ�7��Ԥ��C]�Q߮A���nDc�Дf4�-SN��"Z�6����@G:�9�F��Uw�;=�I/zӇ�)/����� 3��c��F؍ԣ��2��L`��&�M�S��4�3���bv���9��y�gY�b���nY���
V��լa-�X�~���z���V�����e�[�a/���r��������9�INq�3��;�y��\����U�q=��λ�oq�;���y�C����~�S�����y�[��|��#ŗ��o���~F�PK���}p    PK  ў,J               58.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G/�E,��`������JmZܟeG�L��n�*��!uզ��gV���,��Y�$C���'~�\[٬�*� ��0�G.6��s�j�/?t
�\���-�|Uؗ���u�����BY�Քw�~vP���K/���X��0��B3�0�LZ�gh����k���6����*��n{B��	�䯋�يl��tj`���oC����6N4Y�x>���ٍ�m\�3�I��N+�ס���^:��1�4��Ɏ�K��}�:��1���]��/�Ǽ�&�^5�H�l�s��"�<�?��N8��U���W^��^���㏴���o����%.�D��lZ��uɯ+�g;Eo���&q����֕�Z/�OotT�z�����kץ4��s"�����ʟ�z��~l�0����gA�Յ�EV��\��Yw���c��=��������1>�)B?�$|_+��C]y�T�.���if]��0�߈���k�ə�f|�'�9������4���+q���'���r݈�e�{w���o PK�0���  5  PK  ў,J               58.vec�S�Q�}.ڦ�mۼ�m۶�m�I݇��S�t5�5�{��g&s"RN$��{.y�S����N1�8%(I)JS����R�O)*��De�P�jT�Ɵ5�ߨ%צu�G}АF�5NY4��Ҍ洠%�hM�,'ڦ�vr{:БNt�]��Fw��C�I/
�M�ҏ�Y~�(b0C�0�3�����-�a,��&2���Mћ*Oc:3��,f3��Yļ���,d�Y�R��\oEʏ��*V����c=ؘ��Mz��-le���Nv�[o��^y�9�Aq�#�9f�'9�i�8=g�s��y�zA��%.s��\�:7<�}�����.����(�����Oy�s^�W��oy�{>�O|�Kd��Y�f~�?#�PK�1(Fp  �  PK  ў,J               59.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G/�E]E�`��k̙mrX��m-�t=b�����/+Ҷ}���~糕�7f��=tfÃ������:�g�Ny��k#�H��(��k�k�z�i��eBc\e�E��=r��N�7Ya�g}�������;O~9�7cÝ�N,��ta��qs�Mi��-�w��[�dFb��ݾN��,��Xr�ˬ���A��^ve�L\r�ċ<�~6c��E��̒��^�&��/�X~nٯ�g&�x*Y\��``?�p�Ǖɒ�%�j�v]W_ԥـ���>��ڳ;��}��yv�����*����:ʷ��"�U�~	�=��h�q'W�(�������ع֔��A���;C.��`��x��N��=��>�<�} q@�����K��$E�l%��X#�{uiqsi,j��ͷF'˭���)�� ۯ>9fVϙ�w����/*�习��W��u���W/4����	 PK�!��{  �  PK  ў,J               59.vec�eoA�љ�}���]���wwwwww���;$8!��"t8ds2χ���ɆsB�d�_�d)BQ�Q<fB	gIJQ�2�Q�r�O1T�1Tԕ�L�R��Ԡ��j��P[�!��ԣ>hH#����4�9-hI+Z�&eB[�m��Ӂ�t�3]�J�����{ҋzӇ���ʆ��AfC�pF02�0��h=���c<��$&�7%f�T=���`&�����7/��zY�b���e,7�¾�z�Y�Zֱ�lL�&s�������`'�����۫�����9�Q3ǜ�9�INq�3��]���}�K\�
W��un��i�-}�;���y�C�����<�9/x�+^󆷼�=��'>���5��0������C�PK�� �u    PK  ў,J               60.i��g8���W]%�$$ʲ��*�;�D��k"�U�wVAD/�#�Z�`����=��х�n~������9/g����y�����ޭ (ՔT� x�  ޿�[ <���H�@ ))	�=�������=x�f��01҃��l|��,<�`�S1.~aaa�����4����6�#%%�G~���}Z�'�'���v�@E�'�B�����#�»�@�����?����HBJF�/����G@�OH@DDH���� �"z�D@���� �;���|V��ݟGlBVa�d���ѳsp>�
����KH>��������o`hdlbjmckg����������!*:&)9%5-�sF�ׂ¢�d)��S[W����������?08>195=3;7����������=>9=;���su�.< ����#�?.|BBB����}�@EH�D�������C�w$�
��U��B�G4V?��	�����������������#��W<* p:b��o��[8���ӺZ���i��T��hBX�d\��R-Dm8���]��PLͳ%CX����iQ/�$Ufҋ�ńp?�X�BF�r�BB���o-i�x�O�^�dR��n��e�r�/S/"%.�)CG�b�7M*Btl�c�}��k�[��8�1#Z���^��G����cH����0���z���C��_>�4>G>QH��/�w�����7W8}�6��������{~�ޓK�������W��[��*s��΂�X����B%yȲx�A���E��+�Q�π'W?���Ւ���ǴuV쬽�Ή�	��q�']'_���^AIsg��k����������䙰�����#�N�	�L,t՜m�7{yK����QĹ�D��������I��}-���fCd$Lu^��(�P2��M��XW\���X���3h��yL&�/����#<R��?��Ұ>Y����AxsM�?��7���s#��o�.��]\�*y�O_��R)|7�m\�IG��4;r�]D�"�� =��:F��qv��u�}�N� ׶� �7����ӡu"6�K3��]��?���� c	���Iq9_`�����%���IN�Ȁ/ٝ���C �`��/���_#g�W��Xѩͩ��6�%�%�2���sV~��}�{@bZ���<8���[AW���	�M��<E�|��˴��~���)����J�1����!�
��&%��l��j(�2���������%��������<;�Џ3�	��C��%~}��6�Uߪ	�d�I+���kM��V?�a�I�%~Y��]zdkw8x�d�$��"�����LY��x��g��O��FT��G���l����q�U��O�/m������c�TN_�T��ǭ�4U�e�2�-�<<�)��m%�k��&�O(;&oڗ�q�AJ�}Ή*�w��)1�ޜ>g%�����{Z�4��3��O�v;�wb*DK���,m�y���_�2׹�'� Ŀ��æ���Y�}���t�x���/��R����,e��*hu ���|4�G��0
��N+���+���~~�3Rv�g����k�'�����h�V��F7��Q;�xs�F٢N�m�J�K���v j_�μ"f�@*���Ӫզ�F.ѢEZ�Wp6G�n=���WfH����[5.g�<zmG�E"~#�~���"��W6�?���ޒ�s�]TEKg�;��-W����]sʀ '�f1wQD2�`�f��qȵR,�9} �qA��4Ƶ��N%#��Q�Z����7S�$�OOi�j�{�b��#��>	�?�-~_+���ˀ�2?��A�a3�h� 4Zz*+rO�T���牁Z������Ϭǵ�(�@G>�/x'*Y3v����C*^���pA����ӭZga�,����(k�w	��H�y9>��k�ٕ ����`���x�m�ɛr����Z��Q|}q+Ү`�x�����3�}��ꩳ�)��2O/�dO��𙽧B�~ݕN4��9'd#mƥ���l5�9gl}J��QO�"��s��%�vq]�fD��'��0�'���AtI��[��e*؍XEJ�Y}Qr�m�Zg͐a�T�T�e"B�˫�nӓ�j���t�����S�L�	�Q��\�p|,��TI	��=C�Ȏ�#G�8I��Y��;�<��5g���ݖ�*��՘���yziq�I�	�=�q�6�q�Z�l��u�f��ߞ�y}~�pƈ�Y�������QI�l����/�S�ff��C�8��t���Y �h�{>�Z�A�).i���1Z+oms�*��	��\P��ڂ?N�?�]�����a�9���7;ޱ��Y
#Q&� ���~K�1���������R�0ۣM�Ld����f��tt��F��|9�m6:����OZ^i�F�E|`�<d0�Ց7qj���@;���#�ۖ`~,Q.�%�~%kn�>��qSeA�P��MF���o��Eڞڃ�L���ӿ�����b0(޴�ɉY�ѻ9�@�n�S�SjDx����<�T��u�Q�zM�*�֜���ӷQ7���Ed��z�כ=���!d�^׳�!8Q3��8����Y�u)�s�O�Öi,  r�H���xu�M�־Ġ5)|t\��V���h���� 9�Nb�����xJ2��L�`�쏫ƕ�*)0�DE�8QBoٖ`髼�A6�F�ؼ�~�[D%���m��D�|��%r�e��d6����u� �Š��;N$���zrL�D�=k����2�7���ٔ�}������+P�޴�$�`�2 �k57��J�פ}`�n�s�ؾ�a�R_�����o�1�!y�����q���������v�z�-=���^~�l55��� M"�P| ӗO/[��D���&��yT�AX,���P����B������(7����G�;�*Q��4��GB�t;=���x��\9����_�u1;��e�u*YY���r8��]
�%�?U���3�Hw�Z���)���1���ҝR��=`=Nü��D��,>T�����(`��1e�Փ^�l�dXE��&�I��fu���<&WW[3J���.I�ћ+)i˞�A�Q�#R�`�o�+#L��rU"yKe+ �mx��� �����K��
���Sh�f�����Q�ry
�-���OL�ME��5���~�8GZ7%�@I66�$D����|��S��!H��7�J�*�1/��I�٪]����^�����d<�.C%`h.aJ%��<�>���kJD��tZ߶�\�m��?w��2�L���o=YtC+�4����=��<ּt����M/�-�~��x�О��`���e�K$U��c��5��!���/��U�ϝ=g �'{���]��o�w�ϰ�0�e��wfvz�ޏM�+�4˃:>�6���3�U[n���������i�=����չ��nUq���x�����u���V֣,�%�j�Y�$�V��D�Z(����d���)�ܚ������ [����-��l=�uG�ƌ2J;��Wg��W�^=\�n�>�9'� �=G����Lh��<�
Cy��7�뛣��?S����U�ȁ���-T͕^��?��B�=�`<����+��`Ca)����tXt.�X��A�����/mtr�ڀ�,��4��Ş� ��@LH�9�袅�����$�t��M_}I��LVI=�ݴ�|��fP��vI�����h!��U7LݞB���ד�����[��*6�_c[寙}U�=��=� �_��x�S���lp7�ę����钇�m�h�޶�!�k����Z�{�zM����[�4�m�F�����H��*�+
&I?v��?���A:ɈU:A��|�)���(����=������w�W���s�y�ı�K"���x��E�_�_�5�6ʦj�Q_�\b���#����-Xk�z���v�L,��{=*"�U�Y���&���� @�R����H�z�*3�o�4�<�]W ��7@3�)����cߛ���-�� s���I�W�:A����8�R��`�Xr��gp�'�om�~�7c�$��W3UxY{�ȨT�7e����8�y�FK�q�`&!�=!�P��z�@Hzz��F�C"m1���'Q�6>�I����Hd@#�'gc':*\$�[�h�7��yw �v����K���~�����dj�tS�kӕ���R��M�L��{��^A��~(��KӉ%���=�U���}��B�.�`�ڒ�j�c�=C����ťolhz�x�pV�:���>jQ��Ge
$����ks�r�|!��:��A���ئޟ�b�|�[��_�7�ߴAy��?w��biz�{���u�����d��z'g��y.l3��9����� $˙iު�>�sm�F��r7�Tk%�)]��ܼ�G�����j�
����8���ψ[�2���)Ԭ���fb��L�J�!�N m$�Ϝ�=Fq�<���5��X�S(+�7�h����Բ��Q��O	�!<�����i��*�@N�T�M��4��UWDqqO0�H��6�C����Cڙ��v�ຯ�B�/��M���q�&��O� ���x�a�1�^��"�{��vJ��U��d _�{5{�������!~�	��T�i��;�B����Q5��w��nt�JOmj\�� �dS��܂����%���|a{���/�7-�v�L��s�
�i��	,�Y�wL��r���,	M��Բ��]k�`�_Vשs�}_kl��p]��dd��#ٲ!���cԕb��N�����8��)�ٍx�w���ݘZ��e�DNe)A�����p�~��Q��k���j���4�A���ᗊ��6K��!��k�9���_v���r�q9{^�w��0p����dYL���_�Z31n|�z��W��:�pE�o#2�bR|�X��T�|�i%��l���ӧ��vⲯ�F�ƺpl뼳�0*���P��⪲�J@fka'�䊒����3�=�����
el
�彾�y=�S�:sz��>˚�gs�츳Vwm.sP�"ۅ�*��7�W����� �����2��M� j瀁���TUnA�-w<:��#���ƍ\l�-a%�p Y� U�	�~�d<��nz�����s�iB���\�=9�5��{=������l�\���&_M
��c�R:9V��:\�2�D�: ؊X|��<��ĝ7�C+��{[�OqJ�/��wo�,l���� �]X�]�K߲�;�$D�����K���g�cN:�M�=���{)�+u+���&~-����u�ۛ�e~�Bp\+�3�����Vp�q��}^��9wt�-m��U)S�s榞n�����esi`<��Q/7�JŲ��\G����1��*ż�^V���Q1LAr�Ѽ�=���b��1Yel�tX=�-��e�l'�W)�䤋#�Ȳ�L�mc��	���!y/	NVSV�Rg�Zcۦ��S,��C	�ǂ�h��	�g����&^"��]֥ϴ؉a��g���̆�
�,�����V� <�w��GLs5�-�`��'�T�����/��; 2�(�W����h-K��ϰ�>l۾ lzF	-8}�A����O��x� �"���4�����'� �c��q{����g�̴6���s��јJ�ě�eKRy�ր�(s [��&����&L���l�9�K����!��5�0	��D�Ƹ.,�)s2�����zJ)�r��U���A_Е�6�~35qq���N�� {�z]}bpp��Lpu�Ӫ�%���jU���L��
�0<��%�Z7�
\8İ��3t�Q�ɽO�\��+�1����`C5S��l!% �(�LG�FӴ��vP�֛$��C/?3�k��?�/�N9���^M_Y�F�"�^)��8(�EpT�X���v��ڧ�6�uA~X�=����Aw{��\�VV��'�J-�l�zC\���2-H\w�좌wq��mY����Zݻ�Vuž�i�b�G�y�̀+7�ƨ������A�Tf�7t��G	À����5Ŏl�
�{Lg����A��s#e�X��]�ϗ{��w��?}�Z�(����\�W}�h8^�d%�I���5{�k��^����*W�#����9g��
���'�F['b^��#C�8���~�zH�y���s�2����J#o����8�S�R)�ǘ��Л�b�+�XofN]�]s���.5`�׋�����ua�&��ݛ�\
!����uڹ���E�+#f��:���R��·������23�e�'Z�ROWk^'��rVp�������]Oi��UYp}_��m߷1��O�n��B��~V��c�&���M�Ye$���}�{uef:LRm�i����0(��G|��8eʌ��R�n�M*���I�4-3����r�>A�����<7�.�٦����@~���+��w��� ��zZ�	~7��β���"~rZ�O�	������.0�R$R�hq�H����T"�.����!�����#�f���32����:~|���.��EE��,��.�2��n/ǋ�e��ހʑ�2�Ï���촩m��*?��W3
��k(O�W��t$k�zގ���k����P�(��������կ��F�����>/�r�-�R*G�Vg���G��}%��R�h8�E����,*^�m��	J��'6��@~�spi�o�=5��6�Q8���d��1Hn3<i	�Ŭ�R�Վ��Nh!�L������C����f��LBS��~[Bt��u��+E����}�~Bb�в�p%�o���'�(P�~�q���9�݋r�G���W)qAݰ�}I���5�_&c�l]�ڐ���]�e4DT;bM X�gl�w��72k���lY5��n����ד���Y�_@�]��秔�(�PZ�
c��{$�3�7q�*��	�����Z�:K�c7 ��9���3�4nqs�q��P�]��c����'���T.�|3?�As�h�T��5{��o��uZ���M>|��%����>X���1\��33|q�Y�&�j^�ۋ�z�;�B;R���Ù{�n�1����9��@��3C�m�tv0!�#}��h��qI�׍	:�L;[l��R����X�L�@��[5t��/0� ]���)�:b��q��r�\em����ZuW��6R�Ԅ��i2��;yR���զT�89�FhV�IO��&8��_+�>.�4H��]��+O�������3�u�k��zN����^�+olq�7���q�Z ��.�eD{]��{6�-s@���d��y��z<J�$c�����3�#0*(?��f�Hb���b^�5h�BP_�@��y֙�w[_c[�㲺���7�W�ޞd�l[�r�ܜ��Ny[Q�Q��>�a�a4(<���Va����K��:����2ӥ��_�h��K�
�,[��Ts��:��z�l����5�oIJ�u{`*�������Yr�4n�F���O����8�0��jk�(J�^%�]��QA��/.��,=yc��NS�gx��M�ņ����8Y��E�&����к� >y�L�GfJ�n*����	��:����u1��;X���&�����G�����L\6��PT�-��S|��+�#��� �����_C	H����ͻ�O�P]OG�*_�<�e��xX:@@c�#�l:��=���}�2{|��wwz�6���D&���g�̗T�jt��TGo'�E�I��1Jy\�r�]������������W3*�% G3G��x%����V����3*�/s�ғ���Zy�:���u�Vj��^n��W�L{"MdA�'������He��Sb��o���'<�8��|��m�?�ueS���]��B�+���TvJ怈%K
9�5I�*���߶?����r"Iy��}�
}:Z�k������g�PΣ��cC�]����vt,�su�-��.�>�$��a��6`8'wUZӇ4�y���b��<�"8D���A�7f�8$5KnU�15���[,��'�& ����lM��=�����~�_�>�:z�*[���?����a��2/��d�H*��B��I4��7e����_|dsC�@��j=� �Z�.W�˧=�i=*p�	�~M�_F�b�k�}�`�r�}������C�d�V�̘洄:��W���u�����f��J}���l��\./���-�oE���I&�[��H|�R�-�t�ӿ���!\��y���L�T�_˜���2�(�Qz�ޮ4�-���2����#bXU�-�0�OI&B�D�9�	��YP��Lm�B�j�E��ˇw�>[�T�b��pJ�dm�+-���i��݁��.�ղ���H(!J��x�/��~8����ԡF��B�B�@��
�Txo�)uYx��Z��*��[/�b�Z{�;MrƷk�~�ᒠy/?�%��ˍb�l���-�	3�L�"~^�OYI���CME�I�!qv��x}�K� ���]B�PR7B��� xƥ���6˚ci4�I��]�Î����lQc���Jo �\���#�eA�p��s�ڈ�R�#>>��t���E�����&\{�{Rd{��A���L��/��^-1C\�Ho���G�n���'� �S�_�m�f�&&b��8��
�>є�ވ
�u��V��~��[#��[ڡ�`<��M�_m�&�|���cIk:\h�b����6�%�ƅ[���$=n���5������b��g��w��(e}*�}E�
�V�m�kh���T�u�,�g,I	�1���/7������}ړ���rA�}�
e�a����%��ז�v|ْv���4}��7�V�v��.�<޸b����r���o-�ڍ�W����'�'�/���KL_��s:��+��ˢN��|k�c?渋���oPK�[�#  �#  PK  ў,J               61.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G/�E]E�`֖w�'_R�:�������tb����eWt��[u�ш��ZxbHߒu��wLe��=g�W+���U$0DaQ��(��)���A���Z�n�cK�v0:�T��k���ӪSK>T���0�ܴ��K��)��c�<���������40 捍�p+.��v��������iOO��Ӿ`��=r�b`�[�t�<�^7N���x�7d��IƢ�IM��=�#ŜͲ�kq��ے���s<&�7{˕փWU�o3;3G���&����z����l�;��T�r�$����?��S�o�2�>��h���3&~�������i�&�0z�~y����y]��eiv�Uw<Ֆ}���=�D�M�4�e�^���%�;mme�ފK�Z6��-���u�͙{G.lc�Y��׎���
�l�'��Fmrr���	�w�+�s�?4{����[3�bP���W�~� ���>�0>�q��q����K:^,�j:�#���G��GL/Ґ���Snzl��'��W^{�n������O�Un�9�;as}�^U��� PK��%�  :  PK  ў,J               61.vec�e�Q��wv]����������[��;�[��S�/.����3Ynd��W�(H!
S$ˢ���)AIJQ�2���E9���De�P�jT������kQ�:ԥ�i@Ô���&4��iAKZ�:�F�m��ўt���BW�nv�uzҋ���/���b��@=��a(��F��Qv���2��L`"���)Y�T=���`&����o���E,f	KY��+��X�W��5�e�����;6�m�[��6�����bw�b��^���� �8���s�'9�i�p�s�:owA_����U�q��Oܴ��os����>x�#������<�9/x�+^󆷼�=��'>��_"���ߜ���O~E�PKΞ�Cm     PK  ў,J               62.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G/�E]E�`֍��E���9�ɮ���<n)Z���SZ�ZYr��|)Ǥ��˚���!��T����_!�']tu��X�0�G.Vml����������T��.��KBOP���m��{���O��Z{v��;�k羓p�0\~�_�sߞ�~��]ti�X��@o|�뺅�BB�j���U�O��m�k���/�&������22�e�6��1,ݿO�Y���	t�tē�����}��v5K]u���O����|���ڤsizT�K���R����/����6��?y��a���Z��ճ����{�\��}Q����c�<��Vy���W+q�.1���+ހ���=�bN�',n���������fo���g���>)�Y�����A�����2�6��/��d��g�f�����0�Wj{�͗�Z�a��F�)�$�?�2k���&?��=rtK���I�"L�ꗼ�~���>���Ün
��V�@V,XVm�N�jO%�u����<�ٺ�ծ�M��Y��j��-Mk��r��E瘢'�}���м��o PK�2��  @  PK  ў,J               62.vec�e�Q��wv]����������[��;�[��S�/.���a8��F��� ���0E�,�:�Q����)C��,�e9Q^W�"��L�R��v5�5u-jS��ԣ>h�r��]c݄�4�9-hI+Z��h�~mu;�Ӂ�t�3]�
D7��=�Eo�З~�Oy1�n��`�0�ag#S�Qv���2��L`"���}S���zә�Lf1�9�M����,d�Y�R��<�Ǌ,/V�U�fkY�z6�1��Mv�������`'�؝��c�W�c?8�!s��6ǜ�9�INq�3�圻����/r��\�*׸΍�'n��ҷ��]�q�<�ox�|�S�����y�[��|���C_"�׿)�9�����PK@w�4p     PK  ў,J               63.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G/�E]E�`�ǜ}���,�?ey�4?�3�ÃZ��/#?���si���m�ߗ�JzW Rx����K����4�),��`�#3E���8��y}ԍfߙk��l���ҥS�s
���Y=ugZ��oB{.�{���9��?C��/o��V��X��̥�������{������<��I�����?��D�F��{�C湆1��9H<_�<���?~n��y���~W� �E]����]��ylnsU�Wir��Z������̕���V+���at\��v�O��l����_��p�p���Pe˓\��ӽ�J^�������ڗ�����3����v���+�^D.��j	te��K���-;�������>s����Wz|�\�����M��;�ύ�B�rZm��MO$�ra�G�@_���}�+���ŞFV���?���������A�{�l��".e9Y�̖�n�l�����-��_J���tZjׯ���ִnR:�g<l��]Y�>M-w���A����=[f��gz�G`�$��YORs7�}���м��o PK���  >  PK  ў,J               63.vec�c�Q��g^�Mm۶m۶m�mj�Lݤn��O��9Y�ׇ;sfOD��_�+�|
P�Bβ(�,J1�S����4e�dQ6ˉr�<�H%*S��T������kR��ԡ.��O�����4�)�hNZ�*�Fk��F����@G:љ.)/��u���AOzћ>��_ʏ�v�@1�!e��"Fڍң�X�1�	Ld����EL�S��tf0�Y�f���u�yz>X�"���,K�cy�+�JV��5�e�ِ~��,?6��la+���v�+e��n���>�s���0Gl�:�q����9���'�ٝ���%.s��\�;ܰ��oq�;���y�Cwx�|�����%�x����|�#�|�ϑ���_����~F�PK}Y��p     PK  ў,J               64.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G/�E]E�`��	�Re��t�� ���t��D��_2���b�����|�]e[幪����_��w��ƢM]�F���O,�ؾ�����l��m����}ⵠ�ɑr�ʷ꽞�gӻ�������~�M4u9si,j�'6�;�:�4Cs�yu���1۽^�y�0<�vDUZ��G���_7o��}�,�O�֥Y[On�	i�;,qX�K�Ȋ��V�K)4?y���1�^'�Wi���׾FBz]E���o����=p�ɱ�B
�'^���P��u��2Y�T�V���`��������+:�_xo�=��ᦤ��\Ë������-r|y���۫'�bT�I�p���P��������fui�ta��/���r����œ����j$=䖛^u�ފ׭���x}��Nc㿾���[ԥ��,|��[�ӷW̘<���٢	^��^�ї1?d���H�'�WWO��t�՝�/
�[��& PK*���  �  PK  ў,J               64.vec�e�a��gv]����������[����l��O��zd8�ׇ�	��,72W�� y��)�eQ�Y�┠$�(M��gQή��@E*Q�*T���jd)j�ZԦu�G}�0�D#�ƺ	MiFsZВV�N���s��v���Dg��5�nv�uzҋ���/���b��@=��a(��F��Qv���2��L`"�����dS�4�3���b6s��~󲼘���E,f	KY���'VحԫX�ֲ��l`c���6�-le���Nv�;e��n���~p�C�Gm�9�s����4g8˹���.�\�2W��5�s�7ܴ��os����>x�#�<�9/x�+^󆷼�=��'��g��)��M������W�PK9e�m     PK  ў,J               65.i��g4���G�D�#zD���.z'� ����	��d� JD��޻��`����/�ý�9�^g��9kﳟ���ue5e 
* ��o��
 lLL,Ll,,,l\|2|<<|jR"2z =##37���]����OPP�&&%�/�# ���MPppp������������ �F���0P�QЈQ�{���@�o��PP��10��qp��%4� �������a`�������Љ1H���0Iu�������S��A���z��,6�8��T�4/Y��98��ED����UT����F�&��v��N�.>�~���"��?�|��KM�������󵸤����������GsK���޾�����������������������������ۻ{��P h(�S�G.�\���h�X��BA�O1:&��.��)386�|J�7H@���{��Ep��������,������o�% >ʿ�C#� ���������b���!)����9���Q�B��`��H�RH�[L��^����Pg)Ē /�٢���m\���gG�ؘ��Kiqq�	�����u�*�u��&�_XI奫t�2U�O��\��L@_&Dļ�;��Y�Z9]��*���v�e�C[c�-�n�$͆uKJ�c(�p��R��0�����N�E��FHpOܲ����Mv�b]��8S�}�(Q�\\���l;�c�p�/�%?.gm܎*�m����ޮ��?i��N�&�-/�#��gHVX�	���O�� �CNy;�A��&��]
�w��R��Pf-��AkG�u2��N���̒/�4��<��6�j�!�Z)<�o�L�qxS.����F��a�)u@4r���Ф��٧:m������L�WJq�*�'9�OU�<����˜ו�U'���*a`���if7�߹[�"�S����}�ᎿO�EP�����5��ƫ��]�o$�?N:��U��l��<]�H�s\U��z_�� ��`�)�N�AF��������#2ɳ�ʼi�C8�	�t�T���R� �i^{+�5a�&��%��Ґ�����#��s��X[Gϑ�e�V��W��Qu�����I�����堁�!��6?I��-���[>M�:���ϩ��7�[)�	��:G������jN�]�8ڱ�@λ�Z�+%��l]ބ:��q�j�`�pp�d��u�p�����r-�.�K˚����P��ʔr�{��W2�9�o�-b�y��.Xގ&N@w<]�yYζ�N�(�n�cX��������܅�j{0Z��q���S�fߑ�N��S���=��s=�Hws���a	1(�}(o��Z��v�)ů��uaUj���(Мf�|�$�Y"���n�r�q�7U۴��L�+X��Bi{ǎ�kI��/�p�#bV��IE�d�g�����Tr�/��5(kR���[ܠ����m�Q�9��̹g4%A���p�|'hV�/u˙Ͻ���"}#?(��<���{D�A��` .�L������C�K�B6!)�v���L,��^�LG�� x�[K�}ԏo�Mo���
�$P�R�K�� Ҧ��io^<|��՛5�p:�_	LU�؄��Zh����^�ZFI?/ˈTR�4��5�{{�Ú���O_���i1X!'g�	
�Ҟ���WNl~�]U#��۷�y���`���*��S��Tl�yP�k�|�!�]�|�N}Y7it�%�V�C�I��7R�����c�-�gN��2�D�a�	��3 �׌�u�<2,xؗ�D̹h
���{��ڽ�-���
�44�C�ô8Wt��3�M�K�)	f�g��f?\�Q2��VL�q�4:��j%��wM���-K��T�w�Tщ��YQBL,���-=�������y�%�{�Gg�9u3�����'���è�fqF�$��Oul��p�k"�Rz�����,��QE���f�ƙ+���=���c�z3��r�s��8k�!B�t�,j�CG����I#D�z򻓹��΂�޲��
�g;IH��I�[x���٘���~������#r��IѻϷ�Ww`�:C�0��D���<�}�_�G���E�V;8s��܋�9G�}\|H�m+0S�~�޵)����Nvi\�X;�?o%���	)[�FL�4�������gUUK���er��֎@����~8��ۤ3b�)L��=13���/ѧ�e��ui�c�&2%���>���ό��$uC�K��$��X�*���GE��V�j�iy;7�[�҇6v�0�U�iP��Y�b$SI>dJ"�yv�{��R���B̆r��2$^����Zᠨ�<h��Y"6h��=�i��i�%7���܃5Wap���#�ը�)�Z�)
E�E�Uē�2ױ��du�ws҄�{Z��S�
|�J�	琰��[��N�3���Mŋ�J��)�{gۨ�)��wƤ�8/z���r����q��Z�F��YzyI�ʆeF�ɕ�-��vѡ����<ς��_���eK{��۫� �V����|��uoU*�+Q�����n;ܺ�Wc��+.٢/���~�6���L�m��g8B��o$"��AzSyl�`�vI�\�n��yYS�Ǔ\tѸX��4.f[�dlh�q���ĳ�|�f.���v�|98V���I��lo��((��8Q�##Q8�R���tUE{ `DL�R�3%A�aR.Tڮ��K����ŕ�5���n#��O�4U5�G�����9�ț�K[,]d"�����6�:�r�g :��g k��YZEoRA��#��`U�M��M��6=Ѧޚ
Y����S�M�!�Qc�ǲOec=���	gm��ȉ�ڿ"4��f��8 �Oǟu��K����md�k��/=�9�bQ�۝�]�щ�h��~�J��q\_�֖�m�W�Ŀ�v���K�S���t8cˋ�؝ZΜA:\�z`��v)U�5*l�\I@]u��ՠ���tF����s~�y I����U��LQ&�����Gm@��;Fj�z^<�P	�>�L~��W-<B��l
$�������"v����j�9��.g����Ux�z�tiw��O�>�u���{�Q��P.�A�e�^�,�j����2#ԫ@���N<4�e�:V�m��Q�c�ސQ��.�6Wu�u��֔�v�(��۬�7J�<ra��׍(����*����O�õ��4�d�(r�;�YhŹ�t'q�R�#Z�3�����_�K�J̶�v�n���VΕ�+��� �7Z+ѧVf���RAuӯ}U3���fԓ�-^��Y�a���^����!�i�%��0Ơ����{hL��kb��#O���l�O$j^L����_v?�����0�cWмܦӒ�?/�-"�YA�Q�j�r��-�U|^�j�e��9�$�`�d�de��R��_04�u�7[e�6}�=�+l�����w�n_���U���I�<�T�d�v�w�����'�ȷ�6Bx���l��j,�3@�������=�յ��f��n���r��Z�4=���x��ϼ�01�"���x�Z�|͓���5����=3�ͫ4��E�ܶ�]ѽ��|�z��Y���P�b�Z�;"���Q���ebD)!I����wѭ�r�G�����Z5��l�F�2���}�ʑ��q=���mb���b���N�ϴ�PP�H�:Z%F��W������~���lL�r�������J�$�WOJ�A�;�y�YE����r�i�%���dR��'oh)>�6���OtM}����ĺ�j�o|�k75�0i�ͷJ�f�����+�_�J��Z+\W�faj�5H,�+��7��pC�CK�B�Ig���uM��܉�������q����Dㄉ.){z!Y�z�ts��.p>�L�+:(4&��z�;�ٔJ���r�/��Uᥢ��lm��Ҳj���Ҕ��I�)~q%���uo꼑�gg%9
��ܮou[�|7����6a�*[�πu��,g�U�j����ap�mJ�U�7��o���Ȃ��H�m���BR������oE�-�o�d�I�����p�z�ҙ����8��"5������|L���I�R�VfC^J�ja�I[����=L��Q�~�����Zм[o���	��z
B���-��T2���KUF��������z�����vw�����X����BN̜�ɢktZ�.c���<��;4�T�B_��y���s��,{u3�T
���%�E�!���%�ԩ��'�]M)^��6aa��b�;}��^?O��'.�u�ֱk����ǣ�1r�h-A�������Fw��e����⥋A���(�>3������(,���{m@��WC��o��e^k������q~ޣ��;y�c�g��z2>��}�T��,�?X8����Z]a^����dTϽ{H�h����'��"��d�K��YS�i��^A�L�>���.F/Bth�	z�pI��������)�㮷{�}_��T3�OO�:����,-o�F��M+]��tث����l���,����:���g �-�I�-Ѩj�hdYdd�"��g�@���U�3���V����لX����n��Μr��Gݚ�EX�I�Uhxd�M0ʾZ 
���G�S�k*�zD<���q�t�H�զc�K�M9Qj�~�8������o�v#B�8��c	�5�WT.+���3�@K||	�t��u<{�����+�1�{�m���XY�A5��}���~�V�4)
�L~W�5��E�ՙ�p^H�(X�UX��t�~&����|�<�KK�3"8���q)�U#���+�Ѧ�A!vt��d�Z����1�?~SE1��B��
2�i�[�F��k���A]]�Aq[G�a;>_�� ��zM�aݐ��z�}5c|Eq��/L�K#�WG��_~���g���:�X�'ew�j�"�:<���6Rx'R� [a�f�x�	Y��C[�>�r<���1['���V6B����ؗd�L�!�=bx��d`�CLa�hǖ0�Q_��J�Ï�E�F{S:�>��4Z�|�o]����b  ��:�mT�U�ذq8�kA7�8o7k6�j7���n9�e"�Y[.��=�R���h�2�j����F��F�
��8�<�j��Y
 !E. '��>�d�f�ݫ�7�-x���� ��Q�ԁx��_�fl�kB'6����m[�w�'`G�v|�\"6�
d!�fc����.d��������j���^�������?>�P7��.FI���{��d��,�*��6|ǗS��#MNO԰�d�T���Ġ��L���g��O��~(��:�:B����
M��ǳ6U���OG*�����G�f�$pb���v�6� ��C�DZ�Ʉ�/�:	�2����d��P���7�z9{|C���
�Z��tɴ� O��ɽ���>��C���9E������T�[�P<��ɠ={�����O��p��p��j��Rz.����P�W[������S����\~���/���e2\��F�HD��NL9%.~Q/x��}�2e`G}�鉽V�z��v?#�b.��7���΀Kh�����u��aa�˱�{�lb2���Ɛ����H�ɣR����yv7�P��;f��v.��_��K��agy���&6�w4������;[S�{?fܪ�Э"uҝ4��½�S���?4Q$�����DL|C��kE��� e�A�// 	�����C�������(~�F� v�5���oK`;�z$D0P���i	��4-�h���'�lMT�3�n/�V�˄����s{�v �`te�Aܛ�N�^��	9)�W�	 M��3$F���{]' �`BY������W�z��-���74Gz��>��i��O(��~�@V$%��0݆�Z�����"�j��r�aB���9js$ymI����E��WZ?V�{!�s"�ׂ29)e;��I] NM�-���S��~�h��a�H2_f٣��=�CK�p�cb�5�=�9��i��bE��By$�]G�eCN�~.�_�OY�l�]T6�Oz�����~��[A�x���ȳ��7xJ�*��qhmevZ�58�*�)���)O��
�R�Zf�{����O�����Ļ��t(��'-��M	@��;��o)n�cn��l�i����n���Z��X銀q�j|�g�F���8�9E6Q}�m�#1�hbB&�ͧ�H�rN�PFw&��:�M�ٺ�;�_/zct�j�t�L%C�����i5q�)��K��r�Q��e��b���^ky5 ���x����P����H/�ǧ�j�������*�c�lq�8�N�	+��#��.ӎ� �B^ ��`֔?F�m#M�.��^�0�y���K���5���^|�{���"����Fh�8/2Ң���Es��ｌ|�7$L�'��A��3�>]����+�%�1U�@��A ��}% &��U���|�Gҭ�������y~���M�����k6�����ݤ;�N2m������mF����q��vy���YV��J�ǟ�����@O�R��M�c�/�Yu��6��`:�z�V�S8Њ)����00�q$�o�)�ɾ�96�V�y�,�o�d��AQ%=p� j Y����F>�.G^���`�HI����)� ]Ř��u�TSMLf�}tT�΍Nch������JW'�QEU��������,>�$e���T�}!�$��a��,�X�6�ҷ����BY$yVЬ�`����n@}{�"C��Q\��s���(��/Lq�)U4����Wb �m�!"�u�����(�|"
�?�Ή����DƼ���z���V���6�4ԻtÓ�J)_�v�#�L��)����V�G����#9��gY��)�қ7�eN��6��ݞ�
�b�2�&xeE��G%R&M��*�l�_�#�"�^����L�#4�dB���ց4e�T�+��/�[�q�l35_&��ÎT�0`�P����kh��]���2=��'H��/=e�48�4�-m���?0�CX��,0]�ߛ>�]�M�=q&�f��vd��**�^�ǚ6�gS �S,k]���o��#T�4�q��P�{�(ٞҦ/���?5T��G����� ����zȠ2
M�Q���}�F�/��7u.qt	R��^�_��Y�Z����DG����'B,��H��4�� P��1q���&P!�v�Asea"o�O���;75F�Ǚ|�Z4�� hI�F1��L�����Ət�����'?��^U#ZQ��#H�4ƺ�OJAr4"��҅�w�(S�L���g�<F�����G:ۻ�[`���+Η]ҙ+�!s��:y���p1�nh�)X��GW*.q���%�� ByO�kn�,��U���Ȫ���R�ڄ;��#������kpV*�6�q4�vS}䐞	�+n�W����W��kQ�T�1�:4�g}{���-�����a�gB;!���o����ݢＣ�!��M��Q�M9�_2���s�Rg��O�,h~"� ܪ�hN��������?�/Q���)��@Gj�q��V��y��D�o���x�3�N����"V���`�p����=#�n���F.�렿؇R�! @!��G��Gy�M:C�\5�>��ɯ��.��dȇh�сK���<��3@<4S������سG�pa�T"Oo&�Ӄ5O�x]�S<gˈ�0�800��ݍ��e���0�y<L�|���=q̹�+�E����w^~m��w�G�黬}���膋�FP��c��M�6��#>���I�xE�~��6����aI�7�c�1���-F�5G�>}�b�m<n^�XT�|<r��;X�նʘo懦Q+��Ǻ{�������6�[��q{�����Qk��lK\���u�yc!́Zu�v�u����$�ʽ��1��M`�A�Ӣ[�����3`�Rp:F6�1G��w��(��aD�꾇���鮁�8��r,�5WN(G�H0�{��޹��B���cN�Cb�סř(u���o���eL�W���pа8�����H�ӳ�//�;W�t/5&�s19k���5��'��8�*-�5�E�w�*:��cb]։��Ǳ��º��;��yt��ZˤW@�n�KqЩ���J2�U[Y`�h��=�o�[�
�n\uw����RQ�cJ����5�0���낼(7D�:6*�d���p=8
R/��Ӈ�<$g}Kʭ����ӵ�ρπ�WUk�f�~�K[���J�����nɋ�xD�03������>��]v}�1m�y�A���0��q�e��-�EJ��.��Vz��mx\��3 蹱�O��)M�Ѐ.C�l���e�7E���0+I'�B�.˳R�ՅnTO|�0*ɿB��܋�iM2�����hץRY<�*G�B�&���$>���)�}�,��D�WF
&/5P��� Gf]`@V�#�+��\	)���lb�� m�:��D�C>w4��Wٮ:��د�m��(�W�&��u�Zk��"=�x��n|�>�'����#��0I~�@6����>1}��DX��}�� -8����������V�+�C��)��-�?���^ڍ��~�
�_���gF���Nz���Ĳ]���L��Ș�T�ů^; N�I���%�ˡ��=�JΖA/�ug_n` ��,[�_������%C�������MQ�q�)��l��/������58XB6�(��؈����c�� �.��Ԑ����?�֞�����;�x�tM��~�����n$1I�]e���Q��֑^�10g����˼S�$����B0V�=�L�Bu�(4�}��~��"Ψ�</�PK5ר��"  Q#  PK  ў,J               66.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G+�E]E�`��K��J#+T.�<V���h��wc���;W�f��ε�*�5���Қ�E]��D]F���&�:�?�ڹ�
*m��z=�lCڥ{����x��;����5��M9Rbs%���֤]"�W.v	��X��@O|}g�4��eD�c-Z�[{��d�Ѿ�7Xe��O��(��H9����|�Ƚ���;X�3�U~�Ò�������{�b�G���Ó��F�[=�|2>���%���f`&2Xԥ��3/�2�쪊]����v�����7�wJ���QoJ��N��4����>�����g�M\��e�-.P��)��g/�a�_���|޹���k�->���-�b��i���y/���X%�*3^�v���ȣ�܎æ(jǶ��_��Y�ݣ��c���}��'�9��N�%웣����Ƣ	'M'��:V4����؝>���%�3̹v�+?�������~���OWO��ޣ������iK.��=Ð~���i���W+�#_Wj��.�.����IϚ��Wn�9�Ѻj�����[���J���i�=!{����6�������	 PK�T��  M  PK  ў,J               66.vec�e�Q��wn�����������݊���`��J��%��<6���,72O�+�|
Q�"Ͳ(�,N	JR�Ҕ�,�
�(�ET��De�P�jT��]�,E-]�:ԥ�i@C��h�&�)�hNZҊִI��������@G:љ.t�[ʋ�v=tOzћ>�����c�� =�!e��HF���vc�X�1�	Ld������;����`&����2�}��X����,a)�XΊ�;Vfy�J�fkY�z6��Mv�ݷEoe���Nv��=�o��>����9�Q��w��$�8��r�� .�]ԗ���r����f���n�;���y�C�'<��y�K^�7�����G>���%R|����;?�ɯH� PK�*`�m  �  PK  ў,J               67.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G+�E]E�`֓[���d�>3=��*.��ǃ�B���a�޴#2}�Z���$\��Z(�U�$�Ƣ�Q<�����u�%9T�~�w���u<֝�t�ߥ�^�	�^���y�W��%狼�����XnG��<q��y���'٬L��;$U�i2�l���?!����S�o������ޙ�egR��L�����ے�H�m)'��nb��x�Dٯg�yâۯܼ%�s�y��1��O'�����n�}�M��=G�U�.t��-�,�c��c1<���jw���{��I��w�{��k!�H�.,+�����l���&��|��qL�ə{;�ݎy1���YR�Wӣ+�>�}�k�a�Gq�E]�j�D��ߑ#����JS��'�������'�=H��k�������R��|ꡉ��-�}�[�s�DO��
u*�W+�8������2`���wՔ͚��-BK�g���L;�b'�W�^t]}W���E"��:��z�����������o PK+�~�    PK  ў,J               67.vec�c�Q�3mS۶m۶m۶m�M�&u���y�]�d��vn��LD����;�<�)Da�P4ˢ�Y����)CY�dQ>KQA�H%*S��T�:5�j�ՒkS��ԣ>hH�����&rS�ќ���i�r������Ӂ�t�3]�J����z�=�Eo[�1�ҏ�p�@�A�`�0�ag#��c��y,��&2��LIS�1M��f2���a.���g��@^�"���,c9+ҟX���*y5kX�:ֳ��l���-�V����d�ٓ�ث�O��r���(�|���=!���9�Y�q�� .:�|�+\�׹�Mn��m�;�]�q�<��y�S�����y�[��|����_�)��M����O~�;�?PK�P]�q     PK  ў,J               68.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G+�E]EG�(����!�Ǌ'�|�a�������3+s��V����t����)�_)�/��fZ��5�PÝ�G��s�ó>����Z����Kk�r*w�|����0Fg���y��
�����m2Xԥ��3/����j��$���"�+Ξi�K�s��Y�����sS����m=<O���.��g��%��ղ�O�}���c��.+�9褽��9Ua�G�ȯM����וm������(�|��w鹁����wn�����_�dc�+ד������Ȫ����\WZ�l�޳܉�t/���La����evgw6���I6zg�]]|���G�B��|�?����~x�a��������?Wfɤ�N<wr�D���O��i��vD$��qA���x�G�-���W��<�,�콞ʰlW�}6�m��r�g���v�-�P�yݶ�vRg�۫�����o PKR2v  �  PK  ў,J               68.vec�c�\Q��w��S۶m۶m۶m�Iݤn��O�W3�f�OV�Κ�,'2��߹�#��� �R��,���8%(I)JS�Oe��ty*P�JT�
U�fWݮ��I-jS��ԣ>RN4�"��4�)�hNZ�*�Fk��F����@G:љ.)/��u���AOzћ>��������`�0�ag��Fڍң�X�1�	LdR���=��Lc:3��,f3�n����糀�,b1KXʲ�+�g��B�d�Y�Zֱ�v��ؤ7���lc;;��.���n���>�s���0G��Q�{L�'9�i�p�s�w�w�}�K\�
W��unx��v��m�p�{��y�c��g<�/y�k��w�����9R|����o|�?#�PKNNRq    PK  ў,J               69.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G+�E]EG�(���ꉈ�cl�B7�>�#\�~���W��c�<�DC<��<ɴ�$��ߌ�{��XgZ���)d�0���~�?�S�gk��z_:��=o�.S����=r�x�Ѽ��KS"&]zr%�ՀKcQ.l�wK�4R��.�R_��M;v:|�����x�͕�l�=/~:��<��2�����\����W$Ё� ��[���*���3�ͼ�����H6��r=r�}W�%��<&7fI�������f��YV\��^,�b�^����T�r�M�e<����.�|�V����	jk�g(y�����O?��S�S��$�3�Ԫec�t|�M����`�k�O4-;i�H`@�H�+6\�OM��ZkQu�YOTs7�}��=n�o�ëv3�jg�/�8��mމ
��'i.]�h�S��& PK�w��M  �  PK  ў,J               69.vec�e��`�ѧ;;����;,��������	Np���-�4��>���M&"ɉ����!�,�(L��IK�(�KP�R��e)G��$*$QQW�2U�J5�S��v��4j�:ԥ�i@C�8͉&IDS݌洠%�hMڦ�h����t���BW��=�F���y��}�G�݁v��`�0�ag#�}���豌c<��$&3%�����tf0�Y�fs�g7?ɍz!�X�����H���$��jְ�u�g�d��n���6�����b7{�w��>����9�Q��w��$�8��r��\H���]җ��U�q����mwG���y�C�'<��y�K^�7I&�z��=��'>��o�"��i����/~�'�PK���{w    PK  ў,J               70.i��g4�����-$�Q�5F��%�-ѻ�D'�F�h��k��QF���K�^B0�����/�ýw��g�����<�n�n@������ p��n�  $  ��@ ""BbR2RR0�
Fzf&Fz��������y*��+ f攐����"8DDD�$�tddt��!����@E�#��p�p�T8w= ��:�q�; �#pp�x� B"b���zJ .�����û����Q�S?��<ж ����%����v���>b���@D����	�S.naQ1q	IE%eU5u]=}��F�V�6�v���^�>�����?FDFE�Ħ�?���gd"������}�^�����򳻧��?0��������[Y][�������w|r�9;���� ��?���Euυ�������?	Tx����r� ���a�4����]DlB:G������<����&�����E����7���sx@* ��ԛ�ruR�{ē����Fڽ9$���q }����+��z������*m��#�e��dKJ������9��о[��5&��${�ɧ�EP ��#q����Iw5��*z'[�h�mh�ȏ�1s����>�nCz*EJJ����g�����w/645�K-}�| ��%����u��u��֘-\��Z��Ԇ�a� Et�"mY_�׬���E���C�1}8�e�^CIϧ��k,��"y����ﭶT}�|4=s�B怃�C�*��y��I晚6N�}w{�ݫ�%�hjV�v�;'�� ��1��O�z�F�z�ֺߏ��]�W���;��bzT�F�	fۤ}���O��p��;��^ �5��x��g�5T�'��U󢺏/Sh�<�l��IXmT%6^��[�wmz|��&O%��-�Z���~��VgE���2��J���J�k3��µe�)��ymQ�ɣ{�7:�Mw�)��m�hK���㗸Xn�y��<~NVV)O�qG��y_r�~���擃�`On);�J5a����Ư�F���c��W��H�ʚ����r�}��+}5� 5kO��gP��z9��c���b���xX+v=�l����\�t�p�]E�N�O��'�[�H��|��y"n��p��`3NgĨ����	\O}�������<��5kr��
�+���Ջ����%�CC>�s"���?��}��V�=�r�_lp�C�b+6�?�|�3F1e�:3#Cï?�F�5���Z+lVh Ҥ�,��f��\�h��0t���"9�/�I����-�AMI�xD9�GSȓ:qYc	y(o��_`�(�fB�� �7{	Q��T�4��®&'v��߿���f�7�*e�K�N��z_ɰ(�A�5�S��s;��рC�2y :t�'�NR���ݎ��G�]Zc:���*V��������(r��3.q��|���9΁���q�����~�mb�J|�f�I���uA�R�@±�c�
]�`1�^��.�^��^a7�^�����\�����2��r"%/\��W��N��]
���c�W2�R�|uL���<��~E2uD��TZ��rp ��fS鲮��f>{SLU+E��?��oJnp��.���ߵz�� a�%-�������ϐ�X����ֆ��I�g ��k� ��읩�elI#g�-F��pD�G�8dՔZ��EK$�~$D�_��(�u��6<b#�&㵙���StN�E9ʨ�l�?�:�>�ʾ%�2�Pl�M�}u/ ���%P�"v?�����g?����t������p��m��^��:�d�����TJ�����ΧJzm}�{�?)/��q5����9���`���rX�F��S�Q>^�K|9-�?����x6��N�F�=�'�'l�q�� U�^��Y�δS�"�
'�.�5����_��;�;
e�C�9�ؿX�b�;+��Z���dz��&��\��������t��,��oP�|}o+������ǋ�g�WY���220c�����	jQ�i)ɎZ/��x]��V�MG�#�6��Q�K&?�$OK��v�Z��M!�p,Z.�8-�Mm�B���h���V�%Z$9eM{r��NĐ��HTl)X��18�]=�jx��;BQPɍ5Gt�$���FQgCf��<�8ge��*)���ī�%�&�L^�S��C�W[ʄp:���ڐ�Ɠr��0��We���MW�f��һ��/ݢ˟��4j+�Q�EE�a�o5����H�rT�o�1"*�m��.�H��ŷ0����/?�~0g}e�9p�37[�x��UYgPv��LP��u�Ѱײ`�A��2�����G��~��9����Mik���j�_��T����;��p��k=����4���]�1}��p��{�xj�����~~���5cݗ�ԧй��ߦX{�ְ�kw��n��?�M#�$-P�R�GlQxL�D�?�jP5�2$VQ���I�d]3 ݕ����[($��{D���(�u���:����{"���O����"�|�f=� �)3�ܾ�A�3#}��0�]�{O���#��G��t1u{�,@�8j@��0�c�t����^��Q�����7�F&"F�&&�*�?��y�<��`�b��	��l%���Q:蚍�����#��7Q> �3��[e��	*k��#�����Y!�[]�a������8V)o3\���|o"�
¿��$�?ig�g���Y��������we�pRr���O�9��9�n�}��w���;����Rخ��\j��F�.�r&�y��Z�+ӹ'����~/���YaDFپ;��X]؝����R���O��� ��c#��is~U�G�u�&b�_IO�n�V(J�A�}*���n���]�g gaH���	�$�9���TI� 㫂5'��[�}�=���צM;M�]V�dHW������L��711��7|��s�,��~�C��V��إ����Z���=�`Ԡ���B�Ly�����������c��T�v̺fʕL2��j'73�R	�(��f��Ͳ@��x>j3��e�����g#e���}��?ޣ���������7fI��#��e�q���K��C>j�RF3��`ěu�ѝ[.���!K
%�����IHg�ۡ�x�}`���w���߂S���2����?�n�;Һ�ٮ��j��j]OВ )΢D�3ub�@c'�}؝r�9���J���fG`���)��m'��j^�N:��Y�я�:�GD�v�����ñ~�lȗ�sf�/���xj���8�=ƒx!�_�� �:���i�)��]+�q\�֭I��K������P��V�}�'�
�NVV�W݋�Tr���P�v*8*��h)OxuI���C�^6��DW%��T�.�U�@ha#��6<]�"I�v�~�՞�e���3����g��J�.�1� X��.���z��z���fӜ-��i�.���%=�s:S�,fB`�z�du�ڛ��LN��1��`������o��r3������z|:�K��8Z�p��	�O�5l�:��2�Go�Cn�*&Ք=}���+z��qU��+�&T^�e �)*6h�����ul�8TQʝ�K��uyM4�u�����'z��BY�����
x��;���R$�f'�)}AKb�����Vm��h�\?��˩�Dы�Z~������Ͷ���	���r����~<��z�!p����\������ԃ��w X��u��}�:�( ���6|1�3���c�mm�C蹜����qx�]���%�|vJ@���I���?������hP����G������/(��K�t-ɖ�^��iO;s|�xD�l	`.���7}p��ީ��P���=%��s��봰��H�6Х�]<V&-r?��C)�H��i����������`�٨�V??�j��h�|�����S,����S�f�u'���JƯ��m:6�����}6����䧵ā�s���A�����^�B!��@t�IF�6������\�:�g�Y�栤�`��>'��
�MC�[���	���F���A�Ҫd6�"�ϝ�E�p�0e��V"<Tg/JX���5 ���,{=[�Lg���Fz�ֿ�	p����{t��y�Q)W�����f�oڐo%�%���w�W�g�������pF=\"X�V�?��V}$]�+��uvp�ie���!J�q�NRl捣��o6�����ϗ4�azx�I2<�GA�HJ�Ո��&�� ��ߍS4A�+`�|z��*�8S �y��f��Vc[k��݋4�G�=�KL���7����˷���S��|:�gl6�x�ʐYf:�x����4���C΄l<����8�	P�c��&����eO������#oWL�Od1zA�l���XJ�)��;��@_ף�Q�6�R�}�!�:f/�ڷT/�p�D�����(�U�>�4u�H�LR!�l�#tT����6U}fM祭�(�B�a�Ƣ�}��&
�&7j0ㆫ���%����űߧ�hРx�?���LY�x�B��!k�R;e@ӹdhSS���72��z	���|�i�n𹴯#�N_��ׄlê�M�������}�^������_�~�#�pÚ4|������e�Mc�ZXz䵨q��eH��7��Z�y #E�������E+����mI�7�����lq�Ǒ�jQ����[�ywH�!b�~���l2��1wa9[���/��{_�����*�E��"'|x�!����M��oJB������_�E�h��ƶ��^+���1a����nԫ����T�?�3YC��/!w �2>5��b¶84�ȥ�U��t�w觳�������� |vң$�%��o��2+��҄_P��9&�Z��{�k�7��Ϫb��1�6L�����Z��������5�(�dk�Q����u|X������_�
�z�WVȉ����i�2��tǞq�˙��'*$t���𾌔�t�lE��tR�e�N����Y�6��-d@��s�j(M2T{ƃd)c�@���^G#�V���㗿�>��d�ke�oB<��NG�ܶ�Dk̴�o�U�^yb�G��S�t��!�/���~ɞ��y�`6�A!}^$'������|�-�knjn����ɪ��X]�lѢ�x>�'��?�~�|��Gb-8o��0�jt>��)O���O6 ��6w��i]���-��/	؅�ѕ�S5d��|��@��蝒_�PL����; ���Ӕ�-�L��T ���3����V���O7����I*��/H�� Wߌ�y�6��P������DT,W��0�BQ�_X�;����YN�J��R�b�Ju6K~S��1�vi	ǉ���t6iH�f�]��V��7�IӢ��seOwt
����������a�G��h�:G"6�w�ѣ�����ǐ��U����Ďa��"w��b+ۥ+�ҙ@y�z ��$�o�P� x5��ǿ5�a��3i�[�e}Q���Z��?������&z�G24��G1�Lq͐��Fn�g�; f�1��s���i�v��w�YG��d7�꒱t��UD"ΰI#8�g�kũ��gm���e3[;��b�юʛ�ڄ�5Z:|$�����H3��p��ߊ��E_s���I�lL��r}�&�����j��	�.e��2�,��-3�sb=U7�)?�<�hI����ˎ玩�T�v�+a�L���K|4;��9��QWGћo���,��(ϸ��z�mZ/�=�M�TD�2�"��6����jIh��thP�pg��f窓��"�I�Z��ǻzP�sK&�v�&�d�nj���}\d�����R��|+��"t5��e��{�~PM���}�UHި%��n�<�$S�x�/��V�<�+���-��V8�=��?��r�l�Gc�M8;4,���b�E8jL����ՊSH�MP���m���qH�utaQ8��;�%Re�<¥	�F�؟���9���ůt��oVow;�S��}����uZ2�Օ̾W�<;�_29�o��bbn��tۆ�ٱ��{�`��\PS���B��()�F��)�0_w�]U؈&��$�͗Sv�]���Oa���ڽ����>�߾�aaMU��C�v�$�@H�ˋ�p���*���)���:i�\����5�����ۆ�7�2��2r�i����^�<$�_�Ӡ@q��ˀx�ci�,�<U^7���0w �o�K�c��+-W���B`  z�0������XM�:Q��3�I%L�2�2�[�J����|�K��.��% r��D R�,�|VE:� ��HT������'X���cL_�?'ՠ� {
05�x��!'��
� Ƌq��yQ��=���g�H@����C�����˫���>�o;�+��Bo��_���'s�Zc>�/ޥp�SEI�
6�l���S�q�2,�p
��^����\��${j���þG��7�Q��?G�3P�Vʈ���j��x;�aY��)�Z��08���~�7W]+ �7:Q�]�M���uS���as���ـ�L�p��n��[�ƹ�տ�?9���y�&� bv��~͖Oz������UnGR�,7�V.Y?68�&.c6CZ��W�S��M���(�3�W�.���W4��!�r��Fc����m!�
�uek��z���6�]KG�`�g�����.�0��S�6֜\���N��qALz�����z�Q�P�<�m�{��K�I\��Y����u8��V�D
��b���-q��\h8o�7.��1�$ՅY%G�&�W)*>��n���LТU���zS{^R`ۍ:R`�f�!q�]wb��h�[L��B{,#�=��K�U�{ۊ��lm����n�Gn���g�^���
g��9L2S�qfH�e�$�?�KNy�i���U�X+�?eoH�nK��x0d#*X���d�"nCG�TyN,��A�c��n��r�٢�_�.�/2���I�8o�tU~���l?Kn,W_�"���[1<�e���H�KK+*G�����|�m��#�t�x�h/v�ZA��5}��h��2��@�=ӗ�yL�ݔl�ȸ���.��b�vkӮ5�[7�Qw �餷��/���V��b+��*�?<�l��O颎�pP�o�5�u��; ����������t�t}t���XCʀ/�/��$v��Kf�~�2�(�@�HA��eK���$Ca�i�TG�?h��L��&O�4�C�XS�;��I��W!$\?`ka��ۭt�{�h<��Z�_���źZ��+�U��;<}�B��+y�j���+�}䓍OZ���n��Ȅ��ˢ��kTd*n�iW�Kj7����H�p�!F�?�������J�|�P�x���֎�W�����^KI2���dՍ�:��0�o�Y�<�?hv�6�`��*����kf������mz=�0�j̢3�v�b,g��1ک��5��gw���aN�k@cR��L zZ+4b�b{�k��p��%��/	�Iy�J��0�?���=��c�=hޥ i���ى6����"3��WS8u���{ٓ{V��ӼЍ�"� H�UE�k[p�ܮ�O.���8��9Px\�W���	�JQ�����'�d Qy*i�m����*���{��p�u%z/���,J�Eng���!���p�ҏ2WoR�; %H��[C�����?p���J�JGv�U\���bD#Y���㠵����z��+%	�P�h�­?nmyF���[����E��U�1�{��Ƭ%*1��y��XJ5Ο3l�-��5��P��l���.q��@?�積L�^IQ<�G�q��kKq���u�; ҟiS�r;�Z˾��9G��?�o�]X'���4Ѷ��h��aa{ ]Ǝ�g�{v�`X,c�Q����Zw Z�i�S�ȿ�=MV۴o��p�Ǳ��������*��98���	v������{[f�y��q��P�m�#>=�wT��@��T�j�|��SM@�!��"��:�	q��' j82b�X�rkķG7���X��B�3�Ԏ��O�鵻耞��:���f�Uv���Ѹe���e��@�*S�H�ADI�������q�p��g7]���;#�қ�J$��M��=c��2	y�	r�S��,�� J���NT���E:.��L�|���q�����7����~�	��[��ؐ'c'\���@+���ڰt�U��BI5���H:����N��M���7�����-$ jRh���	C�	�W��}j/�*=5smS�A/��Wq|���Se<�&?
[�$~$C>�Nffޏ�@��
mw����v�_cE�!�W����m;�(����X�� J����K�3;�t�G
vz6,�}���'�'f���X������l̈́,Z��'0C���פ-�M�4q�IW�Qߊ*qH>zzW7Mgb�[�W�wu�U7�y[��&:��v�1����}��]��mM�?�X{mB�52�ls|}��z�#z��
�*��6��yԴlCgD��f��p)?�6��	�{ �����H ���b��>�!��B=0�����e�S�"��@���֫ʪ�t(؀7[ū:�#��5L9F�l��*�2q4�2��y�Z
�萢
Ϝ�_]�j�Ŕ�Z�[\���]jw�:ra| J�k��|"^���sv-7O�2��]�u6;�����!�a���=@�#�-^�'=ۑ��W�e�_�Q���F?L,�Ί�/�y�h8~�f�g�{Lkƃ����UY^˄�n�� PKv,_�"  7#  PK  ў,J               71.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G+�E]EG�����?:�&�L��M�c��Se�'�^�u#���%���w�ph��r"����>J�ܺ�pŢ.�@W����b��n�
����!�oՓ�6�����3�ZJYD0?K�8x,j�M�s����W���Ζ��t��<:�������f��SD�IJ]���;>����<ϐ�+\Q�O����uS�V��X4�U$���[_�3k�$e1�K��%��Xg��9vߦ���M��$?6��zd��ľ�.�-,_�]E`�������hMf�`<�g��3�jϖVݺw|���D9�g̒?w�͞~��Ľ~/4�E-�Ґ�}Y��:U;��棘R����~�O5�83m{ٟ�V�[�W}� �J��/��bS�V�qN���+�,g�ږ�
�b��W����?���7WP�qAcQ6|��V�w��t��Sp��Y�ҭs��O*���z��,h�T�9�v�^i.�xQ���U�E����o PK�YQ�  �  PK  ў,J               71.vec�U��P���.����������;wwwHp�C����!���&��iD����=�|䑟�Pʢp�E]�b�%)Ei��ɢl�7���T�"��L�R;�Y��&��M�R��4H9�0�h�ӄ�4�9-hI���=_ݖv���Dg����j���Nzҋ���/�RDs�@1�!e�a�Hs��h�0�q�g�d��,/��Lc:3��,f3��\�;O�gY�b���e�W,�o�^�*V����c=|��6��la+���v���n������ �8l��zT�8'8�)Ns����}��.r��\�*׸�~�s7�-ns����>x�#�<�9/x���+�k��w����_�)��_����~F�PKԕ�"s    PK  ў,J               72.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G+�E]EG��,�Mr����lD�Հ<S�X�O�[�U��MW�z:w��-���2��&�<!�`e�xv][�H�� ���'�H7<٪-ͻ����/�l�����r�߅ROs�����<�v�_�Sve�.
��R�h����gg��sj����jĿ�c�'����^�s^RӼE�Am�����O�{�ݲ��t�^h*��ԥ� ��ۙi�6�D�Kk�O:�����Ŋ�·��>=$Sy���	�����v\�^��;!z��E]�˭'&�vK��s_C�]vo���g���|[��$|�6��>��I;�v'�}�X�`�W���"<Ӟ��'�-Y홧���Һ��+.���=~���i�7���-���+��iҫ7߈?c��^�ҴAs����V�y���K���y�V}�̏}�r\�q����b�}�{>�����G|�KxPx�L�{��j�7]�J=3z�=� PK5�0]�  �  PK  ў,J               72.vec�e�A�ѷwY����������!���C�B�?��əz>�Tg&��D���;��Q�B�H~E�,��┠$�(M�Rή|�tE*Q�*T�թ�r�f����M�R��4�!��{nݔf4�-iEkڤ�hk�N���Dg�Еn)/����=�Eo�З~�g@�h7HfC�pF0�Q�m7F�e��D&1�)��4=��d���\��X����,a)�XΊ�'VڭҫY�Zֱ�ldS�b����mlg;��n���u�c?8�!s���:fw\��$�8��r���o\���/q�+\�׹�M���m}����>x�#�<�9/x�+^{�8���|�#������H����������w�PK���\r    PK  ў,J               73.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G+�E]EG��,Z*�'�^͖qe�F.�I������L��f����k�Y^��pK�v��5�y<�o�?�P��4U$Ёu ����[��ꌰZr~�����_�,�]���Z%޽��{�	�#D�O��nϿпO�%���{rTJ$���Ox�;V焽]4q��_���v\�(���zh��j�u�|�HH�.���wJ�ۯ���|ѭs�汄�zA����	�ނI+����󗖊_��h��x~[�����_g� ��sq�,�E3��OVl�u��R׉�O�N��g�z�����ؾ�U�Wn9�tO:�����?���s>g��r'DO_���A� ~�ug��OV��6<��<)�'��I��^�8&�n[iR��JPYCuށ��SSo2����r�u�Y�@G�O?|qH?�]�{�����k�)�D:��忎����e����[��h�q���v�Z�m�n7oq�Αɷe�3�_Zs��bW�)���:�{��ԲC�R�+�?�y{�6Kv�~�R;�]�w���Nej���,�:�r���DXE=3z�=� PK��^�  C  PK  ў,J               73.vec�c�\Q��缨m۶m۶m��m3u����4��*vWs���w��dOD���'�\�ȧ )D�?Y�+��Q����)CY�rY���De�P�jTO9Qî��Em�P�zԧSn4��ƺ	MiFsZВV�Ny�Ʈ�nG{:БNt�]S~t��{Г^��}�G��b��@=��a(��F��QY�h=���c<��$&��)Y^L�Ә�f2���an�����,d�Y�R��<��Y~�ԫX�ֲ��l`c�b��f���lc;;��.v��q�e�9�Aq�#��Q�c�8'8�)Ns���K���}�K\�
W��un�7�����r��<�!�x�����;z�|����|�#���>G�/��������H� PK��/1o     PK  ў,J               74.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G+�E]EG��,��&^�#lK�Β��8:�0�-*ഛiڨ{d����If�ۮ����߳�o�{آ�/r�)~��}{}���n��z0ui,�7�}/����I%,42>!oa�����Mo|�仕#M�;Evs��K��~n�U57�v.�i��Kc�DG<A��Z�R���������Ƥ4��m��j�I��JB�j.1�+��i?�pR��};)�w�Pz���A�6���I"�/cL��i�q�e���s_������"�߻���=��V$0DaQ�̼��¹�fB碜��l�y������,~����ƫOw������z:���9���ci�+�mc�(�bQ��H�+>\bu��]�OOZ2G�pά'Wj.��\w��F�Y{~��I^]�ݰA�����m�	t�;�����e:�׋z��\�%�:G���I.��?eoR�q9c��,:-�*���38��M6:\��/��ҙ�׿�:�>�Ԕ@W�@#�`ƭ�n��8s�iq��ʃ�������oqi�>�+����+Y �[p�Ә9kw��r�Ϫiǲ��� PK���  ?  PK  ў,J               74.vec���a����u����������V��Nl�[�O��zd8<���Y�9�R�<
R���Ϣ�]1]����)CY�ٕ�RT��De�P�jT�Fʉ�v�tm�P�zԧi�r���m��Ҍ洠%�hM�T �ڵ���@G:љ.t�[ʋ�v=tOzћ>����R��3��c8#�(�7:���2��L`"��̔15ˍiz:3��,f3���Kc~��B��%,e�Y�~�J�Uz5kX�:ֳ��lJYl�ۢ�����`'������>�s���0G8����q}����4g8�9Χ?q��e�p�k\�7}�[�m�p�{��y�c��g<�/y�;}��-�x�>���g_"�W��7���?ܟ���PK,�q     PK  ў,J               75.i��eT�����T�A:��$���B�AR�sha(��!DBZ����f�x���Ɨ�����{���o�u�~�����HEAY��
 ����2@���������������G�����GIBJHFKEOGKEC��������DC�&����'((H�*&)���G@��?MP����p�(��)�_Ѽ���s�E���@%F�<������BA��c`ba���+h"�� ��h@tt4�Y�y 1:�+>RMKLFpR>�l]7���f+�l�/)(�^����s
	�����ɿSPTRV�����704�����wpC=>yzy�����GDFE�$�����Ȅ����W�7465#ZZ�z~���OM����/,.mnm�����_\^]���!��Å ��O����q����0�Å����b4�W|$2���RF�`,2٤��nl&�?�V�8/�7_�������B�������Z�Q�]� l<��Y@w�>�~�>��lj��&=��z8β���VZW��T� 2H�hwW�QO5��j�O︾��S�~cN`#��Ξ��H/u+_���d��v�Y�$A[�d<!r*�e!�ϛL>�4�_�G �1��'�_)^�4�1~`Gⴲ	�o�.ɠ�ٙ�
�k��E�g��� �ظ�����ꯑP_7�t��'�=l���\z����������3�b ��ϗ�6�A+�QBf�C���dh~�^����R��]J�Ȅ�7Ki3Y�,;�l[_h�����R�.��AuA�jN����$rA=�߂�~�چ��J���̀�ڼ��nA&�9�4Cti�jM��/h����hF���b@��3��B��F��3	E�;�#ǎȹ����1�M*}��� ����s���ڋ�M--�wT�V�ޭ��fI�pMGÅlx�����08w槖�C`�㽶'T3��U�ֆ��X~lӰ���}�gA�lg�OI��k6�~���I�Gt��q���g�}eӟ�/���%w4�e��,�m������R��yva[��_��܆�S�K8c�ιg��R,N�<Ɵ��Ƈ<5��B��N�)ز��ZY��i!k�0�<@&�!Y�V�Ws\��.��|K���u��
��f_��A%��d�5�'M�d_��w~)��kP�z�w/����rLR���v��G!H�ě*Ψ�B���v.��U3g���?��}������<��M��߫��aCF��"�/���R�8�bXD^Db�Ò��D�rb��<RkP�M�|��ᭀ�Yu�z�L/*~����`�GΊ㓧uMz݉oǰvl�!��&�q`������z˅��MJ���`/�Z�rb������	WQ� z;e��ħ��-� ��g��P��9��'&rV�$��et�3�����,�E������X�Vky�^���|����.�@jCJ
zE��#t�<����pyz�Qr&�F���/p������G4xD8U(}�������rU!	�s{�x����ߩhz;RMY�e-��E�ru�1������~�{�o��s���~�x��=����zY{o��묖a��'ؘsI����yl�ŷx���%�[`0���A���!���SeR6�NX�i����޶$��⪂��61�C� 4�g_�5������F���")��+�S��)���h��j�3�WbE��E�g�b�DArC*�5|'�sUf��>������HG#,N��n�c�>k\2��p�$�=3H�|�Xf���oQV�qh�u��e���$�d���o��T�նNz���'T������k�pd*�t`�^A���>�~��J��H�*n�){��7�ޮ<q��sO�������"k?�v�P�6��m4��7V� tE��:9q�6c`�g�b�^���2(\QҤ��6����0M�J�F	�v`e��yk��q�/�A�T�b���l3j����l�ӿh������8��$e��(�ܘ,oB��F(���o?�"�M��;i y]��%�1r��>�5w�-���>��sS�˒���6U1D���ªXn����I���L���Δ�@+��;�M��%��yr�H='���'|%���X�v�&!"���)k�$k&���@ÿa�?׆z�~ÉPo��E{�4vĥVȔ�BWs�0W[ߚ�F�DD=Y�g�F�}BfE��!���+�#]y���_�w46���Ħ(P��I�-Jy#$yRp����{:���Sk�ވX�@w�{o}?�K�Q�/h��B^^��|���w����ms�∿2jS�Vˆ�E�"� `?R��x+V��(�^�VU��2q�el�m���F��e۫�3���4���
�q�+�dͼ����iT�6��d�l�me:b�/��g#�Ja'^ݩ�ܫ]j�4^�kK'/�5���!π��G���ڦ ���40Xc]�uv�j��ē$X��7+~��E�LT���R�PU�` �"�:ɵ$2�]E�N���j�K( ��.��>r�@�W���xJR�
L�x6��٤g�G4����9">(���F��k���v*�4lC�p�^$@�wx�t��k�ib:�Ć���G�f�=�ϝ��
|��P�"�f����6�w������ ��(&}3�w��yza�g߄E=(�Fj��S�c�:��ޟI��)��	|���j��m��.̿+��p�4�1������U�{t2gz��q�&.\"��r���[�P޷��&t[	��WT�m�I��+���s��?�,��l3�_	���k�mKkk���|*R0�������/��������l%h+o�x�$bV��4]+6�Qt�;�}N-l�q[��*{�k��/�'
�7���-t{��|JtY��'Ў�?�����L.w����I�g��H�k1]x-Bi6_cY��=����j��}
]c[0�[ ��Z����;.��j�ƙ��]�턅��GJ��@'��y���&�'�ɩ��V��f7BqU��n_�N^�;[J
�r���d�o︻f��e\�F�ۘ�mC��r(�G8c�P���-,N[�j3��ـED�����s�/[w�C�exJ@r8����
R�0���{��O+��g�H��aW���~�ۛ�U�Af=<���SJ��;R
��z����y��Q� ��ù�x�sM��c~M�Qf+�O jU(XlN�hJ���W�*��$@�hp�ZA�TE#��C.K�K4��Q���.���Z�����{�$���\�弜�ܥ�uCW"�j�S��1�$��U����O�kN��E��'?ړ��f��44�z7�S�&��&=���P�͝L��婙Z�N���2?5����.'e�����(�y�dZH�ż�h2S�t�(;)g�RG�?웗��AqW��@ ���b�{��gȲr��0ʄS�j������Q���/A��Ӽ�昧�^V�?� �K�)�^Wd֨�E��)6uMkh$�v!���ȩ霿���7.�"q#4i~��";+��D%c=��ǟ7�)&���ֆEE�+�#L�����O('��F�U\�ҽD�����$��2�;YS�K>���i��0�����eR�%׌�P����q���7']�s5߻�q��k&E��Ol��}��(n����g0I�2�����4Q�:�T[$�B���~9c���E 	��F�'�e� ���͍�/�p+Yv�1bg������b��ͱ|��U��X�A������۩��A]ss�����"��A଄+���lu ۷z.
;�(P/�`+�8߫�V�j�gY�w�ـ\��A>����/j�����>C�&�=ܖL���[��x�5j�/f�Ct���(jJ�@����ii�."�hi�Ǝh�Cy�﫣nUmYcg[���J�Dón��Tf�Z/��;nU�C�e'��C�{W���%��L/}���D�X����4�(�Y( IH�}2!�i�T�C:��&om��*�fܲV��0^��/5��ȧ��Vg獵}$AFC���XD�&��Mv3�ꁷ�R����lg&U��>�O����=��`8��QުL��j
vҐ`N�:E�)NJ\��֞�Ms(��*(h˪���N�# 4��2]2�w�-P\�����{���%��V��3�2�#�����h���`�ո�{��!����م�E"AqFv@�.��M��D9�o��5r��d�q��=��&A���Ϥ�Z�c"̫�n1;����Ⱥ�E���	
�OX2E
^���F0�'rFK�C�k~u����R���^sx��,�������%'��K�1@���+\F���t]��{���>,7����?�\S��U��>���QN��:Ϛ��Zi�(K�Q��S&k`�g�=
L��7D������ef�o�a�[�?Ce����2=�9�B1w1� ���Ku��u��k������M��rM�;�'�81l������Dف�f��y�!��;/�}�uݪ��!��$�$�
��F��t������G�]Cv��������}ئB�*�߉|{ل�cvKDMi�ny��QN�v��?j:��>蕳��7d��I^�ӻ<���4H?���'E�ȯI1�}��0i۩��S�����K�����W�ք�<�n̵��S%u��eUb��ue��M��;V�˺����ܵ�
�կ���N��n�ؖ�����٧�W�Ȳ���-�rg>���ҁ�c�:���ް�1P�kR��I22 �t!|�O��5R����8��������9���;e�ހ:����B{��ak��nu쮊��H]�ܒ�q$lB�
59���-��o�f�<��JGD�\��w������W[�?I���_>@�WB�G6tMu���\>1���U�	�V�6�krJ���, �i�/X���$�x_h�O��W.s��� ����Y]�s�g ~��'��8���m8�#�B��Q���ZXᕒuq�ZB#�H���d~q����O��(�ڳ�c�-[iU�'�|mvm����92r��"y��Lȹ�ç����F�_N��#Ȼ����
�Fa�:�"�����o���=_P8��
�3B{V]H8�m_ky��X/ʯ4c�F�5CMjAY~��g��.�G�`�q�O8-�O���	lx��Ҕ5J��応?&�/�V_�����u�@Gx���������J��h��C� Fo=�~6����&�m?ᑽ��杅�T���;�^�;X;�J�$�qp��\�$Ǆ�ِ��tD?M��C�(%�7ѧ1�iSg����Rˆ��ƃ\�p��*�I�:`���49���9�x�1f�(֝�����J���E��6���b���.\z������3<6�T��y�����j���I�9�|������Yj�h�8 c�i4/	��B�Sj�/B�?��zy�}������D�3���Ӈk�0���.�ͻ9��B�2�~j?�%���bgmW��R�ISgW<�oރՏx*�>d���V����i����,#L��Xo�I�?N��6�d�ԫi��K�f:l�Dx��H.]�W�YZ�`�ߥ�����c�����pu�.n9��'��H�[�ye����o���B#$Pr���l��đ�cy����e���L_X�%`L��
M����O[m�3 �7��0�����L+��B����6a���ϩ������EO�&�~eVZ߹^*����l�U�R����H}n�Q����>'�S���t�5π���.d��RL�{����.M�Q�|W�]ii}Uu��0������5��oh�1��R 6�H�a������&��w1��ڋ�j��2ؿ2���Z\U��4�͵�]j�jJg���H�t{�}��c>U��C�ԏ���TZ� �a�UW	O�D�K�nO"�F�������J��-c��g�Av ��RC>�C'酌����oJU��]UNa�$MC�����S�\���-v�r�a&z����K�g@0G�58�����ء�T�� Ut���y�Ч9�j}�ɐ�%Te	2��}8��`a�e���BD�Ԯ����ݣ忑.�d3IX|��b0w_n��:���]���q8^!ݎU�L�L�-@�MF�*����c����P� ��]�e�#�h>�]���U����8�����e�]ԩxY'���'d�hL�=ZK�����C�>z X;�~U-a�<e��6\1,0�N�����*�j��ȅ��hOJ�=�򺆑�c�;�?��I��:_H���N��-�s�Xk@H��_{�͌���л�Gp�B3������O#7P���aD�JF~���6�/�������s��U����Վ;��k/.��I��d��'k���FA�e�:�bS�h��U2/j�J:�J�>����L�z~�����)����|>Ί^E�MmB6#��;��҆�x�b�]����`+Z����
\���C|íꎘr�Iws�<7�����������ܰ���YtL�̖!�dD�e����D|���TԔA�����c��WIA����0��斸�$��0�1?^/?YW�&p�J�%��La���M5[�э!Uv2z�Ǒ�_��;��co;�����G�������������v$ko��ڪ<��}5�Ui.�����o��M�{2���=���F�ilɣi�����{X�_�������~*�O�����s"���n�y
	(��1�Y�}��x2ʿ�i=��˳Iѭ�[
��c�=5�ywA��t�x��4�Sۈd���,@��	�}�qb]U2��q�(��;Q{����j� }J?�?[H��6t�Sٞ����ב`J5�� hhk'�� ��`��}��$�V�Vz��������uQ�ׂI� ��lgƃ�ŅLS��40��(bj�A�g��ː��g�1�I(�����\��t�Z�1l�Y��m|�-�܆?���n�ʛ�� .�I� � l\�q!2���%t	��8�ͷ��
j��SC�����G���q�0g���Z�����R5>eƏ�cf?��>�e����i�:�P,�P���m:w� FAiO=qV���?؜����c��(|@<C5�U�YF) J�=��>�zB/<q�ǉX��/.Nw]�,j���j�`��l�tu�ؤ��X�"CJYa��~�$���jK[t)�����JO�,�@	���2�/B� �#�\+]7�!Y4�rФ�]�$�a��
*unN���[���'��ux�_�ך�VR	�c�:_�^����=4���O�g#)���xҺx;��Վp�oR��
��r�G�����,�����Z�d��g4�Z��3�~����H�*u~/ӼC��C�8 �%ɾ/�y랮F~F!�
�]��h޴��&ʗ�مmF?Tb;o�J�&tj����jH`PZj(g͛*>���i���ߜ��0��l�Cy����S�F0�s�~ۈ����v\`��5 ���X�0�r�h~�O����Rhw/�gH���	�(�ZA�j���J]��dV%d����?��6�����A90"V�U�8(���2���������f8����e����`a�`�=��`�J]��P?��m��qcݫ�ͻjS��0'��y)�91�^>{Ă%Dɨ�O��a��ᗉ�	X��%�Nj�|���ѩ���j�"��b�y�#&�
�$e��j��T@[�����^�SQ� &g/5����[Fߋ�2�%�;C�q:k٨�=V�����1������o��_�)I�;���4�/�6$���7	1�DT�Tv%�����F��{����o��S��׌�#|E������s�u���Q�l���t�,�2��*���{����I�>�/���̇��)v�Fߝ
*7y�#v���pw��n��\m�c�M�ɞ��(l�п=�]�R~|q�dd�rv	��G�;=����!ǣ��%�9�Kx�Q9p=�!Ծ�BJ��
��Id�Д^aq2�S��D�Y�1[�� �u�#��&�T�P��臍��!xN_g����
Ny4�`�W�}�)�z�#��:z��B$|j���ɉmsf�����ӲO�!*9�I�f�S6x���G���Qf>��;�S}!�����遼��[��{��]in\��ݗOv����7���T����(Z�ϕe���S@bJկ��_ɔ�J:�3�J��1]b.��JT���ؾ<4��NJN�=4X��@g�k��aӖ���B�[��5.m��J��NP��u�*W��8�B�h+{��-�P
�����"D���bK�������C�O���̢���`���}���sA�
̗	�Ӈz\㣺���BVˑ�F������g�~
��_�Ϩ9~������9/��[J������ c��wDm�K�
e6T�}�=R;u='Q^U��^�k�j�%�u|��N|(�;����
�}���<����>����UFw�h�[ee��e��56�E�E��~ЍJ�LX㤭�\?�5�?��Hu]&�]���.]�Yץ�E"�2�=�v���P�t]�Zt�	8F�.Zi����JDic!}:��u�d:M�I���&�e�D�����/("�	mz�?��F�ۉ�
�.���*������g �*!�]]�X�iZ��������~�ì]$]�ޝ�+Aę��0q}��e�`?0 �����/Xwq����$Z(�����a�m��́�8�=>x0v��iC��)�D�bvm\Ɣ�t9�����PK�U0�"  9#  PK  ў,J               76.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G+�E]EG��,����-x����l��ضk�J�>�Z���H�u����^O�����*<�<���^W� �@W:b��e>+���`W^g��4{�.վ���'Y5�gx��s��_7���h:����K�Il�b'ߞ���D�\O��=�3��Jr4:.��fT��Z���J���^.sr=��h�#�@bw]qG9�H"dW���	��1)���-�u���8�H�u/+��un�Kڱ� �b��}�]W�|Ns&y
�iאP��x�+����E�x<���A�Ў����\���D碫��Ƣ\ت6���`)������r�j�n����n�)V�0>_�΃���`��?��4M8ԥ��	����}p���cM>so[�>�`��_��Ʊ���b��f�?e�W�������/�૓/��t�Jf��*�~:��6��]�?��h�c�ε'�J,�p����o��m3Wh�|:v>�@�_��s׾�ū����{r�f���.��8�+/u����l!����eO�U��a�Z���zϲ<��K#;�w����=)f��m����� PKED�o�  B  PK  ў,J               76.vec�e�Q��wn���������ݭ��]`�؊�J��%��<6�3Y��r�#�B�E�(fW\��$�(M�R��v�u%*S��T�:5��r��]m]��ԣ>hH#��h�E4��hNZҊִ�mʋv����@G:љ.t��S~���{ћ>������b��`=��c8#�(F���7V�c<��$&3��)b��t=���b6s��<�?� ˏ�z�Y�R����L�c��j����c=��&6�,��m����v����a��>�~p�C�G9�
��	}�S��g9�y.x��v��e�p�k\�7��m�p�{��y�c��g<�/y���k����|�#�����/�������?����_��PKSh�cn  �  PK  ў,J               77.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G+�E]EG��L�m
��Z�>yg��l��lߧ�{�"���bni��m������\I��5iǒ�&��&��:��K�g]Z�9���1[�[�S^do��)寳~�63��U�BO�߳�R2+ߧ��sm\k�d��������g=T��S�#9��Q@�.��I�mb����jW7�2�6SD�I�����t]E�D]pᒪ9��V*
VV~6X�g[���������̺>��*��Bg9�PW��Wz��q�E�u�sW��әxh��/�����Ϡh�0)��n��bK����d�==u/_֙I+qG	��N\�pa�ڴ�谤I����e�v,?8��D%<yͭ�r�^ld�;�wg��g�՞5]$R��V$ЃPg�����Ք���N����OZ�tr�ǽ増_�jر�2ʬwO���g�?��8��l�M���u���%ƻ)���Ȯ]�5�������7Pm��iA�5_�/��m�#+wl�<��!U�gP�i����iK�5�(�Bnc�}t�H���[�%�3����5��EV��Yv}T�Q햙��ߗ*<�n��oֵc�Y��o PK��H<�  I  PK  ў,J               77.vec�e�Q��wn�����z�����.��.�[lE�?���aq���e���!�<�)BQ�Q�0�v%u)JS����<�hW)KQYW�*ըNjR��)'������O҈�4�iʍf��\��%�hM�Ҏ�)/:�uԝ�L�ҍ���gʏ^v�u
�K?�3��J���c8#�(F3�=�f��x&0�ILf
S��}��w���,f3���c>ҟX���"��%,e�Y�JV٭�[�ײ��l`#��̖��V�mz;;��.v������<�Aq�#��Sa��;�Oq�3������7.�]�W��5�s����6w��=��<�1Ox�3�󂗼�u�o�oy�{>�O|�KV_#ŷ�������ߑ�PK,Om  �  PK  ў,J               78.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G+�E]EG��̮���%�Z9>�������.]�{�1r�%�s�B��k�/�3x&��
�{-Yת�*㢫�2�Ƣj`��,�I�J����ew��-�}2����/!����v�z��=��0Ù���㘭7�ui,SXԥ��3'=3��ٳ�w_�m�SO��\w��ooWM�&{��6uS�[��V@ږ��ߦ��()��p�D�a��F��<����k�;�W�w���<��'�<s���������i��45��:����r+����Tٳ��dE+�h��%5~�~;m����[�x{�*r�N��~i�%�}�o����s/��3���zc_t��w|>����I�,��wj�K]��40��|����r}�:��,>q<��_�qû��N�ۮ��Όl�?�S���g6���(��Yԥɣ����}˗-W�v���3*>���驷���<��[���z�uJ\O4��Z5�<=ȝ/�R��E�yK�4ML�ը�Y��Y�Rt�����5[�]nM��4�Ⱥ����&��WZ�pQ���V��{��܉��B�g
Ϭ��W���%�ʀ��ӘƩ����!��Nڽ;&Wk��bX���S=�+��I������+�f];�����M PKH�[>-  s  PK  ў,J               78.vec҅�A�o�wgwwww������]���
�`����O�1>�<|�����Y��<r�S@1�S��EY��"J�e(K9�S��T��^�,EU�թAMjQ�:�MyQO��܀�4�1MhJ3��\��ޖr+Zӆ���=��st��Еnt�=�Eo�>z}�~ҟd��"����3���b4c�8���&���d�0�iLg��ff1K���2��,`!���X��b���e,g+Y�j�譵�:y=��&6���lKYl��!�d���^���:�C�G9�qNp2�)����r��\�"���sż�5�s����6w��=��<�1Ox�3�󂗼�5o��[����G>�/|�}��S��O�_�o�D�PK���l  �  PK  ў,J               79.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G+�E]EG�(�3f;{���]����7�>x�;��{�GcqE���?�%��mq���/�P������2���m��cXV�>iqLzi��^�3=8�t��8p��L�0_���f�+P�+*f#�"�E]80��kO����iKO��v�	gϿ��Y�>m�զ���'^��~��@f[���K�g,Y3�;[]�7x����MϜ��~����Ņ��#�m�<��L�Ƣ���"������R�W=��v�EkT5y�g�z|��-��Q;Z��O��zPǙ���u���'�/4�v��H̢.M����K�L�5�������_�i���Bڿ����U��>;��3���9K����1�?W.]�h�-�t����Eq�sRU�~	���p��Ӱ-韖_�"�tƤ�v���Vg�g�]�'��ʎ�rK���;訲����a)�f,�j���G��>�ؓSk�
ш䅢'�+��|X��n��E��R~|0��s]�~�߬kǲ���	 PKӵ˰�    PK  ў,J               79.vec��Aл/����n}vwwwwwww�-�b+b�)y�G��|3w؍Ȳ���K��(�(^�E�,��\�Ҕ�,�(O*�U�RT��P�jT�5�E�u�WW�G}АF4�	MSn4�k.��%�hM�Ҏ�)/:�GG���BW�ѝ����[�C}�G0�A)b��y(��F2�ьIY�5�8y<��$&3��L��t��Lf1�9�e�Y���B�.����,c9+X�*��Y~��ײ��l`#����m��&og;��n���}��~��r���(�8ΉT'�wJ>��r��\�"��wY�|�k\�7��m�p�{��y�c��g<�/y�k�d9�����|�#������E��)��O￬���PKY��'o     PK  ў,J               80.i��UT@��� ���%A�7����F�����!H��ݝ����y�����xNժ���ڧ^^6 �d�e H�  ҿxYH0��1��0100��0_���`c��R���(�)(���ԴltL���s����D���9�y���6)..)���^� ��Hb�l$Z 2>
>�K/ �o�hH�-��2
*:&�+�	��H((Ȩ(hh������� T|4Nq�7�&�N�\~�9�t5�D��ܦ��X��IH�����Yxx�>�JJI����+hji����|13���jeuqus�������������_PXT\RZ[W�����������>0845=3;7�����gk{gwo������������.$ 
������2**
*����������FÉN ��a����P"6����[�/����+b0�&��������������o�% 
ҿ�C�@ ��e�3b�]����m�2�G&�#{c�y�C)����Y�ÒJڴ_yj3�<�S�'�	��lߠ▔sT�����<#��no՗��[��#.kޘ�n�@�Į����c��C��4�On2�x�y0�Z�2�i*'�& �lM�>R��&Q�>��nHE>M�P^��pT�F?�M ���=TI�u�`����14׋A�4d����x+��(˼�U6�l+R�p��.��蜳�ny�V�
%���"��/�k�xKn����;��l�,Ǌ���[��,�t}X�*�X����C��Z3�N�^�6�|z.3�A�?����D5�����-����:tv\��T>ߠW�-A���RNS����|9@|&�bP��;0�M��h9�T��i#	v�%[��ʴ^y����D����܍����K�Q+�Ѕ+_-5(�	=׹F�(���pօ%`�Yz��hw����^���gIJ��ץ�E�3�H꿄��
��{;�v��&�e֩�Z=��e�[�ydh�ѭ���&��F�A�1� �nk$���U��<_iU�j�AbE��<@����n� �ս��K��yU�#���Y1�0ަ�Ր��X�h�n�0U��y���4��K�ʆ�Z�����WذH��ۃ7�l��G0��.��X�Թ��]���Y!Cʄ���Tq�Op�O��~�JA�yO�q���ͣϠ�!�K���|�<X�WC�zeo�41���&��D^I:ԃ�������$����h%�'����0T3_����Q�<����k�*��l.�$�R��<�mo4�3+~��u�p=V���};�ZB��#�B�;�1ث�,�5���T/���Y"J2��� ���H��p�!~��� `y9��s�l�>}�8�{L�N-���@X;0:�%m���Cu"z(ݽ��l��"�BO���MY����G7:��o/ N?ĔB��i��a�Y�ɉ̎>{��4G�Y��S�̕A|��m��T�X�Ws���#��ݝ�ߎe�������*��X�?Ɖ�����􌓲�:^��y�̯˭=�5��U��W^y�#5���-�U�"٫n��Em��
�k(2@Ո�j��w�>�	�։X�d�p`=�g,}h�=�>�O���.�<�����Io>PU\��ضZ�qQqb����E��������u׮���ju@����mb�v��SbD9��8�j@�K�h9j)����ӏ�*e��F3��g�w�m%�dbe'DG�g��w�){�LC�v~�!��S��n��/�{�7�M��3�B�jy+��}�-�T�+v$���x:���7��M��-��:�)[�'��o��ҳ�-T�щj)&~l �����H�IJ�PWѮ��n�!���~�p���]e�\/$�p�j�}��uO�Ӝ�97x�z���.Q�����b@�V��|SF�#��7>���f���#���PL�|+{���f�^(1��9P;�Ƕ&@������έ*.�����b-��1�ЊY���r�Oh����`r϶<2'��J,;
!-h���A�)��ڜ}�%��=:<D��4������gfY&g�F�B�>mT�'�:���w�g~���l�i�����Da\�wLi�W���� �O�~�;_������h�)<jZ-��ŧ��ȡF<��kE1�)��=��~��]ᖙ�x��+���d���`��)�d�Uk�Z�wvZOs�Zϐ�R?Cf?]��r,Ν0qۈ(V��q-�=�V��C�o���h7W�:�.:_���޴�~��$��v6?�f��ΐ$ޤ���wi�o)���%�7%�1�V��s�~ȣ�`�G����(a��~N͑�!8-�%��i��b�:�8o�g�S�Y3�Z҅���@����o��z��(E��J�tDF��.vX#I��aF�ͭXc�.��)v�z��d�vБь:Y>&&*b�f�Ld�Yo��Y�2�ª��������a%"��D�@�cO���������g��bl���njh3��{8��ݜq𴚻�p�%�>KAe��7�q'C�}?Y��l�48z�Y�*��m����>ϸ+�(�(<���7��3b�=����6���HѳH�P��2U����i��S�z�An�U��l���Ov'm���5���`F�,-ՀO
	����h�X1����g?`�Ĵ.o��;�����EMbWˋ��yVV�n�K�t���b��РT;:���T��q�V�?j���c�m�
0f�!wJ[��K�˼��V���R�o�\��<�v�[��T�Oj���3�݊joϼ�y����{A���ߏE�[��%�pyn��m�QL�U�na�P�[�CtL� 1
B�'M�b�͵9�/��ޚ4w������O�h�����?睗4�q��e�4��ͩ��(q��~7�0�MM-���2;����X��L��Vb�y޿Q6�i^s"�^ ږs�����(1�����?up��ҀH\d�h����]]�,W:ĬP��C�Q�k`!��c�a�?�����b1�Ϫf� �(���8oU�C{&�ñƩnӎM����'�	*уrM�STpS������P���=�h*6d�v^�Iɰ�,N��=���o�����kޅ�g3�_Cu潁���4˷U�e�5�*#��JM�ʌ�W�Zi��- 4�蘐<����l��i:��`��n�9C��&(�gYЄ����2�@jG�u�~�meNb�d�ގ��j�3KK���sp�>��c�F� n��=�T��s�wō�(ZN;L^��P�Y�M��+��ѹ���_!^p\�䳄`�]�\�3閆�߆?5VϪ�Tq}��.�z{"'㐢<���X!bʟ��2�B�9xb���h�M6�^��k�~�4������.���&W���!,���f��`�z�Ul%u�����J[.mn�.ֹ-�
4W���F����Eu�K�;!��*�})	ܾ�	WÈK}��n�[B�[�����jm����5g�檂6�~���6ۚ �r��3����$�$>_܂�l��C�����غʜ�ԜϼD�Z���eW������g6������R�Ό��Q%�z@�Q��d�mi4#O<���s9.�r&^��;=�C�i[����.�e�?4
�C�|,j����k��K�Q��.�2��3V�k�N��1tJ�W1_�|0+���[0UG�!����z�&r���0D:�?����t]N�ɫ�V������	5��2��6Iw�Y�c=���|��2�ɜ��o�����a�*�O��#��
V��2:6������+tnL#?=E'��j�o��VR�U��'zn�E/�a�Pm�]�ӌ��CZ��v8������R��0X�Ն�v���Ġ���-o�>l$r̛�E�Y^�
M-�d5/֘��'ߍ��UPw��G��SC�)��z�RI��떉��X��`��|�݂L�z�5�@�Em*�^���|��௴Qj�g`��a���[��;���{�4k��$�h���x�
��d�,�=�gm��c��U���& ���>��L���mXB�C��s�C	�]ZR��`���8{��]��yj�g� �/�/B-����f��0�o��*��e5�ҟ6
|cټ���8��hF0i�c�yG~���S}���C�S�Zx<�f��F��H��v�Ym��D��I������!�N6��dp��})�UN�� ,�����dI.b�qh���~�
�k�>�t����]��=��5Ǵ��i��\�#�~%FX����xP1^��.3�D���.�"H��ʮ�bh�)$-���d߂�Y� E�qm2��엣��y<��^��W{l�3i�}���x\�D���~��"`A��m���i$c+�h��`�@��ϵ�����U��þ2;�#�ïx����� ���g��2h����x�?����^F��������Ʋ~����J"��/r�~^�T̓dب���z��-ƍ^u�U�'��D�8��s%/���zԎձ�� ||�6>>�
c�?� �*�~�s���p�Lq�Ю��2�y�:d�,��L��0�����L��� $~NL�L[��ŝ���(�T�[}D�� �� ;_�;G���M�3G���	Y�JP��J	Hҙ_QV�sc���*������;N!gIE4!��bS0�X�W�X.ř�7=
?k��۷���F�#��	��-F�+��&�Mh|#d��=^�;hi*�tr�,Ѿ�)�D�|@B�-UB�X����v�g������)J=����<8�F��R��t=n� !�.�`ˤʘ�S@�^�E�0]����]�b+�w����1��9*�4tw�S{jE����%���=Wa������]�.d�Z�2�8��L�h�ھ���tR��m�W���;��r��&�~�wF�X�Y�����ހuf�����R�ыcs��#�v3IuS:�����T 2?"�}�ˌ,�����twB9X�<H�
���7Y�̰�j�{U{�^m^�@�;����w	����s��\�lQqk�yI�ɳ�F/n��~�����Tŵ]�X��;��o�c�wo�����3����.�8V7�]gM|�b�k>��ſ'WL��0E�+HXH����� ��P@��\�?\zԻ���I�Q�ZkLA�b�+\Ύ�>)����_$����NO6��1����{o�v/55E���K���ic\+�x�TOן6�l
�&~~��P�ż�y���%�a�5��wb��/˪��~��}L������%�_N��_�B�{�0���.�¨���giN?�ZJ���J{��0��i�ݭD��$Jyj�G^i\oU��*��U�ɫz'k���3f:�S�`6�Y,UԿ�� P�V6���+� [�F)º�k��*�7Nl����3���.}9�0A�:,�ɶ�d_�T[��������_ا��MS��U����үD��mG+��\eI7���H�wY��sp���K���M��z`	�����0�{�:bAا�:�����\�� l�z=��zFQN,r2�n��v�ͪ���HƌW�B��!��.��UjXG��g,����٥
�pyŽ_�iQ�_(_骉���_-�q���?���f�l�ʌQ�P߀��R���0]H���q���;��r�b~�;󾁧��� 2ίV�>����D��۫����� ����ڨLz�=�|ބ(���Kq5��	/ M!tƙ��8-U#���|�؎������9�=^iKz����۳l������u0F3wH�G��'P�x�"Ǳ�`�����Kq����W����^As����t�U����o��+�uֽE'�p������/�ٸzZU��N#ER������>�	R�V!t����Q�*�.�Ŗ�q�bYGz���2�>4r����8� : �5��-�=���;/��9��A�.L������d5�+mW�F�G��]��x�.�<�H���Œ��ؼ��3��P�M붻�L���{���o�%52�� bl�a�R{=�Lظ[`��R��?wf�DG��kt�zt��cmbHt蟇,��g #�;F���7<��	WK�z��I�������������I5e��q��0�A�t���Y�$�6�Yl�]��ۉ��T�v��E��|\�{�De%lU�C��
��B<�83������	L0�R���z}���/��r8��[w��ϝ��/Si�{+���B�@��,�Y�+U(2�ӆ.�/�"|����b5��O|���LUb��d��ΠQ��S*m��ć!��٢"g{j���J�U��'e�>Ԥ!�u2ҁ�-w��GVW*�됅>���@�8���́J��ߍa"��u�qF� |��.��{v���˂�4��	�䚠��Gq �����I���*���c�u-Cc���Z�VJ��1hS��*'мUw���oe��Oy���:�Rǡk���2Xn�n{�)!�!W�1�xF����<L�;��?%ՠE��K,�GNY	S��m�S\z�aB���2��26��x�Z�%���w+4i�rø���E�*_KJb���([(�9���I%!�2ڐ���d���X~�D���YNxf(���-?I���-o>�BJxNj0�"�I���r|O�4���&f��6% HR�uo��VOYi�'�)�������;2�{-��G���Y��NJ�R!r�8��>�"P��Hw�q]bj���ـ�6�it��`"�]�  i,>^{�#�L3�M0/@>�߇��d��mUW� H�\�k��+u��4�v}{�	���E+��P�WǏ�_�]b_��ie��o�^�7��z�e�FW���(<Y=Z����]lHKh+�4�ѝg�����N`�`�]�epV/��ҷ����9:�X�9NwH�M��@s9��Dp�1G�u��<N��JE�2D�G$�*ؘP]\�W�W0튝\��w�l*�g/3�G��/ d���\�3e�g����µ�����׃nO
���u�t���O�v1}nЕ-H�f��,�6I�3��i�ï�ֈ��̱�?���,fܐ�3��h��Pf���UX�ԡl�T'J%@���A&1N/��#�E�G8�����w/NH"GҎ��/�/�<�6x��'1glkmS��)����Q�j-6�$e[k�^o+�5���m��{5���$E�%G�2K�^�@����[� �ޙ*g�����<&l��iX:ė�)�Ǔ�'ܫ��jnA�x��5�9��U�ʝq�*�(��ڟ�Em;��+T�W�.���_a@��X�u���Ch�'
�m���w�Rr����:"�Dt �t��Α�(��쓫đ�Pw A�o��<ƽ6v�̭e:ߗ��E��Y�|4�X[֛�+(��Y�m�OF, |3s��Q>"N�(�t� V�	y��Xʤ5hq�6{t���0.��� ��j��޳�3E9v��aqc�FI��Gp�,�3�,B�{27D|�KV��=��b���|�r�@�x����Ns���M��G�����.j�p���**�5��T�P�_m� �Ku��-Ҋ��Z�y�G��(�SN���6��<�|?h��*�Žc����y���(�ä� ׼��
�PVfbd?���W����� \.���e��k"o
�D����K��|w�b��A��Jbth��)0nnK�RCi�
��|_s� ?�?���H�jUe}PR+��f�=�����p���=�X%�n�e�E'��ϋp#�t��g|jNظ\�=��@��85�,%��1���m��/R��#��"8 4ڮ���1��A�j
ʓ�|>�W�dw�M�;���C�zn�Te�o(V�A����Z���Ƀ߯�D^����(������+E�|�3Au�oH�b'��}sfq�Ucr]쮲�\?��@����.c��;�g�z~UrZ�b���&�S��ALƫ.��<V�.�?�����>�i7����\�p�:9 (�s΋cI�|[���j�!.����N�TZJ6�˕��0
G'�h�g�%�|n%G�n9��=<]^W��i_l.Gi2�]e�J���e�{�A#��5d݁��Qk��6]�����C\�����󠈑���[�7Nk����#���z��>��_
�>k˼/��ZC�ddU7�!3�B�m��M̦����?$iw?��B�4+^[}�a���S|c|D��1fl�E0�� �^�F���$O��h�#%���=*GA��'�mMC���z���Joݍ�E�֘��AG��z��kr/�`%�g���cx���d^��Y7�Z#��c��U֨7�>~�<?nC�b&�y��ΨT�3�C�jJ���Dھ����D.��c�m1��d��j��-�`;7�4��*��z�*߰b=������{�\�ߕ!!�G3��~�~t#�G��E;5�4ݦ���,�p�Gi�۷o=��l2�9��PU���� ��Q%Z��7�E(�k��V$�WV���l�2�J�1˲���v,����~J$Y�Pv��xG򩞦S5o�k�uW�h������uB������~�17ʼU��Զ�,�Y�?�\�6��1^��e��-�F�3�_˪�uE����s_�b���:����N��w(�o�me�ՏB:�o#L�����y��O�
�"`���$��Y( �ik߅=S������0_��s7�2�?�+��*�����BI�C�GP�pF�3�;�)����%�+>�ʵ?������P�Y�������=�-���r���#���m�\܂�˗��PK���"  5#  PK  ў,J               81.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G-�EK]EG�(�f��V2��yw�������%Ζ��X�Jb�O����>��J�"�����45���z̧��Q�|��b�羏��g��f�
ҩHar��*�8�2&���n�"�/�i�-V9յ��Q��EO�_��/��,��qٻ���y�\��g� y��_��x���/�ب��dƢ���a՛|�;|bp�F��۳G;f�����lY��)Yi*�S��O�� z������\�QLw���3,�����]}0�������|۟6�{��g���Zlxe��m�v~!2��eOl֮��*{:$�հU$Ё�5�x�8;xV����ͯn��r�v�����u��]������@��n���O.L�h��s�UD�{����uǵV_������Zk��
;7���n��c�z�s��Ow�8�����v��/��>�^�tS�6������WJE��D]��M�>y������Ag�/���t��_�4�n�Nλ���[-�o��ܯ��5�~���7PK�@��    PK  ў,J               81.vec��Q��;�����ݭkwwwwww7��-�b+b�)Y�G���.o2"����C.�ȣ0E(J��,�g��.I)JS����<R��te�P�jT�5��r�vQGץ�i@Cј&)7���f�9-hI+Zӆ��Ky��\ݑNt�]�Fwz�n�,'z���Ӈ���?h�A���0�ag#��1�s����&2��La��i���g0�Y�fs����'d��P/b1KX�2�����Vey�Z�a-�X�6��͞w���z���Nv��=�5�����8�!s���x*��;�Oq�3����E3�����U�q������]�q�<�������<�9/x�+^��o�oy�{>�O|���k���R|��p�S�ҿ#�PK!�Ds     PK  ў,J               82.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G-�EK]EG��L���vF��T�x���O�WX��Gk��ݺnm��
������q|{ i�;�4u%qi,j�'65�82?�F]@㿽�_ץ�Z}��J���7���c�X6�]٫Kc�¢.<��썱ّ�.!y2�����~�>ꭩ��WE&�f��1�HV���(�=�F��G���͜���UX�G��o����;���V�y���i�$O�E�/��?����ui�l�oʢ��JQ�V0ui,����G�n���=�$��3M�g�cU�7�=��3�z3@����ڨ��g��\� |e��H0>��}����FǸ'ObP�)`l�׷t����A�N|b*����mg��J~U,���@W�V�@V<X��Ôc��'3�̿)��s���9�^�	g:\k4Uz�����E�~����Gef�\���U$�D��7��+c/U֫o�������<;{��y}�}O�z��i���Y��j����1��ۧ;TZc4�VJ�-���"�U�f\���u���������yϏzi�{��g�%C$�Է�~￶2�����7PK��i�  9  PK  ў,J               82.vec�e�Q�=�����������]��]�
�؊������a���93'"����G>�Q�B�ȟ,�f��\����)CYʥ,�g)*��De�P�jT�Fʋ�YD-�6u�K=�Ӏ�4J����5��Ҍ洠%�hM����z���t�#��L��-Et��!����C_�џ��$fC�pF0�Q��v�1�X�1�	Ld���75ˋi�tf0�Y�fs��~��,�,b1KX�2��Bo��*y5kX�:ֳ��l��lna+���v�����g�+�c?8�!s���w��|����4g8�9��\0/r��\�*׸�nr����.��σ,?��x��������|����|�#���ϑ�KJ����n~��?#�PK�+�>r  �  PK  ў,J               83.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G-�E]EG�����_	�p��gǣ�}���*�n*���v�^f؄�L�w	�S˖9O~��7cÝ��.��ta�#f\��9K��]|�O��}�zw������!�/��VI)YJ��2qi,j����'M8�\ �&�����_�r�j�fo��{�j�N����-���)�V�U��R2�h�fsz��3[������:�I�[#�wƿ�v�uz��I�������E��3��gH�v���O,gƢ��@W\�d�֋�C2]��*rݑ��+\Z��9v���|�Uq�"��v�+=��g	㝋��y���g ���_W�5�d�-��!q\m�c��űi�3u�-�I{xg���<?i���Y�������\t��X�ŀ߽�~ɬ��"�������o��V�nz�b��=?�B���n��h�!R��RWpVմ��&;�L��U"�(J���F�_�n��]=۷����I����Sߋ��$3�����K-ٽ^���PŲ_][R��\	tu\�+m�\{{I���sZs��0=k�>����6�d�,C%�Է���mm�ӏ��o PKC?�@�  A  PK  ў,J               83.vec҅�Q�3/���������.��.l[l�V��)�]���6�΅�Ȳ���K��0E(�7�bYA�KP�R��e)G����JT�
U�FujPS�VQ[�C]�Q�4��Sn4�}M�f4�-iEk��6�G;��r:҉�t�+��"z���{ћ>����@����0�ag#�h��dy1V�x&0�ILf
S����ty3��l�0�y�O�cA��E,f	KY�rV�Ro��jykY�z6��Ml��bne���Nv��=)���O��r���(ǜyܾ�INq�3��繠sѼ�e�p�k\�7��m�p�{����xd>�	Oy�s^�W:��7�����G>�ٿ�%R|-������?�_��PK�2^p  �  PK  ў,J               84.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G-�E]EG��,]&9_���5DzU�.u�]�̙j�Zz���83#��2���'������l����T�}K���ftA��xn��k��7�X�m?q���_�*��'^}��Y]ʩu/��^��J�;��Y����ȋ;��}�mZ���ȸ��uF�#���V�����*2M$Е.1�vF�ft1K�\6Η?å�X�������j�����je<<O7�g=V����"�;_lk'E&M�^�=��'����~G/�u��*]����[4�\����A���??z���.��lta��/�:_tk����7)֎猢��xɗbz3[��޲K?�4T�$���\�9^rƖs�5ӝ�D�+{�:��I�Bڟ�+<���sZ��M��c�"�r�2�g�P7c]Ⱥs��i���ۮt�� ���z7���]��y�Ӄ��R�m��>�^�ݽs�-����~-��j�o�h��vIۮw�UT����MW�2:s�*z����eŢdѣ�d�?��\��nŧ�N��O�3�|���5��M|����_W���O�m!Δ��'�zC�"W��#��i�{�^�^_4]_�T��$YW��㯫k;���� PK��  r  PK  ў,J               84.vec��UA��ܻ�ֵ;���\������l�[������G�;�2s`&"I���!K9�Q��L���D��(J[��,�ȧ<�H�4��4��U�FujP�ZԦ�^]�֓�O҈�4�i��fz�����iC[��>�E��r':Ӆ�t�;=虦�K��܇B�ҏ�` ��78��y(��F2�ьI#�&y1N�&2��La*���'3��b6s��<� ���H^�����`%��$V뭑ײ��l`#������6�����b7{�k�}z����9�Q�qܿ��;)��s�<�9�s��\�2W��5�s����6w��=��I&��y�S����;|m��-�x�>����H�kџ�f~����ʿ"�PK@9�Bv  �  PK  ў,J               85.i��eTP��n�RPd��ni�����S)��K��))A�:���x}�u���p����{���o�������ݯ �)�*pp �p�P �����Q����3��R�=}d~��������������7/����0�KBF\P�OHX�?ApHHH���((�1=��}'����++ ��� ��O�����������C� ..>>�?k�?; ���晀!����`8���M���^w�]��3����#���\Ϲy�ED��%$^+*)��������ٿu�8�s���������STtLl\JjZzFfVvNѷ�Ҳ�ʺ���M�-���{z����S��ٹ���5���&zk{�����������?\8 <����#�?.\||<|��p��~��5>�3B9"ZV�pb:yham	�������Cv�U�����7��X������\ r<���G NԳ���rt�)=���n�(����P��q�U��tB��|�3�iT�,�5>��2�j(nɠ�2%��\%
D7��p�^�C)���J_�Op-���un��=��
8�c�X���9 ��2�~y�NX/�hWp�0O��I*1%ɛy�X�k�Y� -D�bu_��m�@�' U�Y��߿L���6ų���~��H����8ى@�1w���0�mF4�6����iF^v,��8fq?!�W��ɬq���r����E�Z�Rz�1=��S��&���߻�u^a73�ڒ���PҖ�k��i�*(zC��ȧ}M~|��^"��1L���W)(��;����E&�Y�T�ج_:�eR�l�l>Q��:�)vZ��>�6Ӡ�a�
4� v�j(�kT.������Z�� �>�N�,g w_��@�,�f���h�kl�n�#��t(+��Ϙ�j�.�����R�m��)�[��K����2	lfO����F9�}�r������l�n��[;h�̟����%��W�1��T���VG��a�7>nX\���!�]O�!��)	?��8T��|\�f"5|\�̕�|C:9ɥ]��=F ��]�H�8'�Q�&���U����嶜_D�$/V���wqW��c��o�{��mD_�~����/�kHO~{U	���*㌱^�_	�iK �4���[�zj ����p��|"q���8�h	g��ս��Q����T��]�W��0f�#8��CD�*^~)�L<,��;�L��B��S�_	z!B�N�na���Ӓ=N;��y��o��X+bq�<<��Yc���=|�v�;ڨ�/�\�*m��>�L7Z���d �R��7�<�45��GQ*{�庱����D~�2h��ױ+Rw�0I{����PI����H,襙���%Ҹ�y���@?b���[����<d��u�q��ȷ&9�F��';m����Kh�K�������8{�j���,L�	�!��I�� �Wv0C�%^l�r�B��6c��R�4�)�����s���&g���|2�)�3S������{��!��5��.���:/u��TV�*�=b��<��T�Iyb;������7�0~��M��s��l�	��b�p�#z�>"�p!�����~Iv�W�5e�U�����2����ig�,{��=Z�V��iP��'xo�C�3��Q婌Sua�4�g"�V9X���ֈ�9#���iJ�9�4�t���!j*��������F��<*3ClZ.*���A���_�p�I6��U��'vevz���ǜ���9��/m߀�Kn��CI,��S,+w��N�Ua�vC	F�}; z���[/Ζۧ�}ܜ ~r�M����؎	��諩j��4�� �n7^�GN�����h�O�Eb{1�g�p8����}�R�� j�t
��cMd���>�����>��ҘU�y,�aXr���,+�,�{��o;����=�T	���`��Y���	-��T�S�:�M"	�{��Lne�r<O��+�o�X;�z&�;����[)�T����;G��T�������(붴u{�Ytp�+R]�Pi�Q�WP-�(��~hWs^�D�i��#
>È�>��d�vr�U`>��vXu�]ᣳ6?7�fS�$���!Ô��|�E4��]����˕~(/*�ܹן	J
 L�$��6�y�H����a����d>�~5vН�N�Pk)�۹�h�!�T�z*��F:L��?:�D��=p��
7�%���e���_yz��U�[M	�1��
�!�gXl*���l�+��{�@>��cF����I鮩����]��궯�{A9�=�o%|.l����*/�K�FE/YK�'��'B�F�1ݒ ��(Ԗ��%�w�_	T/Y��kb��*��G73�-5��f�n�g�Ő�˻�!eZ�9��@Ù�g����繸t	D^q�.�
"C��Oge/�criI[F�gzx���G�A���rv�E�"/:����G?b����Gӏ�?�A�Z�8�iL�^����͎�+�;z��G�|s8a�(�=�&��$�Q���f͍���Z��+�u�vS�nNE���ӿ���ݜ�Z	8Snq@,�:t�ԡ�����^��K�_p�Y��
�~F��%!�'P�I���L4,�>~�_�c(�ZE>2iUz�ʫ�1��3�}й�5�����8�:��uZ]o��I�zA=o�~ow{y�Sr��X�j�]B_�W:j`O�h*�Z�g�n4���Lb5%>��[�~���`%���Rm�"��H�f�ҩb����������w�/�*��K���`�Ϊ}'�`��Yͨ�J�?T)��ʁ	�p�C�Ǭ�mm����U��]ѫ#�E�y��	O�cS���2��5泶G�]��]��=��2�s0֩�;'nh������ʜ���~�8<��X�(��yG�$��8R/vlQc~��-��˸Q�@W%�X{0�T2����c�bq ~�ܰx&�G\��N��wq�"bP&6q��-2�g�R�/w�P3 ���m�i��7�Э"yq�e���˅!�tYu���gO�_4�J����:>�w��f~��ل�d���P���:���~M���;4y��S���]�Ȟ�
�>�m�I�1\��c�Ou�Ƀ�o{(ܷ��H����ӝ�'4�QD�"/�ɐOԮ/K󲢬p�I�t�e���cͫ�_^�z�u��
e�Јq�6W�����@���3�K����-&�m�����6^S�?\����&�4n�_~�x=t�ú�~����c!4Cֆ�*�6�ƶȊڂR�ls}�����V�f�C��peUu�WT1��}R��[��ߚ�O�d�T�dļc]3�(?}W�%��Y�}x��|%gu�&�����Ǳ�V���ڍ�g�`�K��'R_*�c��!�k���DZ2uю]�����]m���r'4~���=o,-��?�BЊ_ݖ��ɛ��UgJX��N�cj�'a��W��7.н�����O6�d�'1���BV���YUI��k��*��=��f3��F�s��Q{�ݾE��5�5)� 4�`��(�0.aH����L��'AO/��qTu ��qk��j@c@u��Z�����!����S�!^M�'�K8�zT=�t5m(�;T��g�E� ��ZTߑʨT���7[�VC�ս��F��+���)�Ɗ�@q��L��:.!
��J]{����@�~�{��خ�r�=@+(��Hq�/҃���q��7u��g��j��"*�=�y�����=R��y� ÁE��ťX&�x�~��l�T�= 6�kT�K˲�����^k(R=��Y��,�·����Bd�qvY�-�!g�m������w����e�]���mjZ� �W���1^R7���Ӈ\��$L��`n�nK�I�f���,�U�gJO���7� �����E.�<Z�#���\e@�~��٪�eϒ���&����Z�ے{ =-��@�SV2���p,([�X8�B(���n�)��Tu��A]O��o �\Yc��#��p��i��J��D�jT���RXI�0�#����2Q�X��S��B{�d�O�Gj�2���Z�/Շ� ��]�k*���?I����P��`��m#(�n����T�v�4���x�_�P+k�}@a�7OHO�cF>5�{s5E���a���Y����ǲ�7��F{��xr�C�T ��^��o���O*�t�3�*A����
�����"��KX"F^L�,=���:^�Ѻ�bۦ�K��a���M��g�!��k�9���؀�4�p'Ȅ\Q�Bd*�m-������0^��ff��j �V�v!�a���7��:o�����ʯ������Y��������ͅ�ȭC�1�#>�:O?����Y:QFiO��L���ʀR���״�M��\iJ}��í���c����f4�;%�l�9���mA}5���J�($"���n�r�k>z#�2c�\`��P�&�����e���<�|p����������+�������Ǿ��&��-B1v[�Vwϑ�+�r��3�,F���/ �1z74��gݞ�S�L��u������B+�Ԡ�Ĳ��2�3�g�� �IQ��];��)~�9vbd8M�A��*U��fY�Q�?�
�g���j��*���B3Yj��s���k�q{�L�����ر5�w̾@▚ϟ�z��"X��㶂���Ax�@��V[s��·)7�ѯ��
0ԇ��{@U��Sx��4���1�J�/����@jE'Ww`����+�U������.)ˤ�����ۿ"pp	����ۿc��l	��H�ϊ�%$jYt�̪W�<^Y�VP�xw���ޱ���B����p�����5
��o�CM@@l����FP���KS�E�Sph��)���,���(��%��n;L� ���=J���{��$bZSD�6l�
�� �dM��B}U��T��{�=��L������f��1�����o��C�#��|T\���s~��j�(~�փ#q�X`��+(F��U�啕�:�@�����wB��Ks#x�j����46�M(������^I}U�]UY���G�J��gU���N)�O��,UO�����/��*C5�RM��2x�<���3m���z�##�v�O�������,�a.u�be�ѻ�t��M��$m���R���x�s8�F	�ò|�S��#.Χm�U��؍u!�x<x|��		����I�7��N��ՍW�����ؕǽU��3!d�9Ԅ�Q�:��P��!5?RZ*|Y:C�H�Tj�wy㦨A�#@��i[��&L4� }����%�6�B�c�2K�p��`m�;�0:�ͷ"SfK��tGT��w@��8A��a'_$Z�VY�-������'��F���t��U�ٴsw\�~da㻍{�o)Q��?����dנ�}��/��mS_��ۏ��d�������L��!�/b,������s� �qg� ���2�A� ��RˋC�����<�����L�X�;�欻���F	��B��U��!d&>�TuN�{@�V��WǙ����7��uJ��d�EqJ�9��������i����bVH~,�� ����U7s���E�ޣ×@�u���F�a��=׹��)� �'��HS��E�nr�q��x�|�^n`*�~�E�,1��������|o�{]������K�k�}:ݙukc�򢇶P6�}6�8�����e!"�~��v��PV)�(�Z>y�p�`�=`K�,x�t3��i�]z-?�����7?�o`{�=Py^4�4?�$\_�.�"�N��8u�.?���'"���<x���lNb���7���K�VS��@�];uZ�}���n^M_�_tr"=�&�;d�8�t}�O�^o0�a���w>-��y��%>��)Zl�X����Mq��D"���v�5�/1��s5K壂!:q	�
�"���g?⥠""�v�C嬍�����\Ӭ�ᆓ�O�$� gǱ
�d��o]R����N�9�&U⡿&,�]#�,3p7oP��<%��VB�|�\�3���3�`K�w�o�w:@t}H �4 J�:Î�O�\}ڲm�;�����/Td�:	�2t�< ����.t����.5�ҮK`Y�WDO��=�����j����Z��4��WH��R�ے�rg����YFF�
��$�nA�[C��~�K�rO������L�g�ƚ���1a7������~(�����F��F��f4�+%���ں�_�s�r)�����֨���_�N[<��	;N�Zϥ�wh3�z��~毑�G�Pgv�� t����,�t3eBF��!I��a:iΛ�,��%Xq�<�l\S����I�ɻ�!kI��_���-�!��x�e�qR%֚�J�O��+/4���Һ4��3)�� ����g �攼�i�w��PZ+��c��k"Ԙ����uG��!��;5�V�'^f�$��0#��wa��:͉���u�/���+e����T'���)��|{�ZPΐh������C��Q������z�^�9&|z���3��a�H
9ZdZRu`r+]˃.�:[���ƶ&���mJ!9 mbï����`���FU��F|\ݾy�ޝ/GbNUa#h��T(#u�S����Þ�����ͺRL�{@A_�w�yFLeRyնN�t:�
�'Ե���k ���'��-""K��*~�x�~�͕�_�Ყ	����Ü�xZr����.`�Hv����Y�ΌXH�yL#��J޲��[8ڍ�sg�����I^�t��� ��1�y�jL՚�$6 i�#���V!��$�ƕjO#CR�p�D"X��I���#b���|�`����ϦVJ����:�3����67���ߚw|5}H�b��������S��֭���7�LG��%�mE��Cn�3Y~\�����3����4�smO�
����K��#�C����a�@o�`z��2o6|����#�>�x�rՃ�5 �֨W
,ԕ��{@b�sK����O�ƪ!�i�ϼZ� \�<}���׾,	o�cZ̬���֩�Mz��M$��\�0ܲ��r�ݔY0�C��j�J$��'�1��ٷSH��G>�f����՚,(�U�d`g�M5N`���3����h�x^tx#,�+
~k�����+�z��<L[S����9Áel��4_��Z��猶<ΡwK ��G���3�u�u}Z�"�rR� ��s��h���T�����d�1?BLp�S�݆�kK6c3m���v�ņ���<�-��������!�HӘ sy�j1�ƹ�0ʝ��a�޷��ݰ�p��qhi���d'��Z(}��t��x����^�a���Z�e�$��z�B�U'�k�,<=�X!)J�'�t��l���t����z>V��p1�::��MG�i��&��}�{*r�g�8u7\F�$��~�.�����l����%!���7��w�USv}V	�V����|���e� o]p���L��������E��ѿ~g���l	�+�禵2��gS�']�ݕ�T��'"j���Q ,��4�Q���	��ӂU���!+��b��V��XN���n��JC��O�D�КS��2
���p�j2�A��!�#����Riߕ+
M�h��<C"��H�UG�k3��%jz^�͔��&YV����a����!��P̈�[���͏���VxL��PI��X��EF���4Ð�C��L��hs�!���ӫ��X?��`�&J��Iyy�]/o��;Ϝ񶪲� v��O���q���G4�{�pV}u�gݹN��0�藲���/~iV᝖��><_�2��c�3��m4-�]I��y�N ��M���!�5i{#ЉC�z�<��|��i�!�Y�6M[��ha	�c�G�� Wp���<l,N������t
��ߒM:ы3�����孑DH7ƐmhVH�ǃ� @�v�6��m��+ovhT�e����fY����F	�+�|�*b&֥s��x!��^�C������40~�S�'WS�੺V�v���*d��c�t��Ш�����_D4�[��?��B�	m'���f��"�[ح�`7F�Cu��E ���媦Q(�5��:�f`���"�ۏ%�d���{�@���_Ga�ݰfBb�x'T���i�\�~.p� DuJ2W����t;�P�@�tF�+���X�ټA�E[��5r6���-c�'a�����O�o��u�&���P�3�-Dn
P�?����몰�Е'r:�R37Po�����
�,l��D��N��}����d�:vn�'1XЗ���m��?��v��CM�|���Q��*y1Uҳ!���z�E�>�N�l�4c}�,��1	(�i��7}�o,�;���ɨ=�my��xYV6��NnK�ӦӇCA���x��Ӂ��X�@�e��.��+'����b��b�8���U�Z��W�������C��= lZ������sH����4>㽣ϥMoKh������*0#����e���1-�595���� �}�>:�z�7MJfF���/�G()-���a8����LB.�v5T`ڦ�I�^�Nĩ��zH�e���܄l��|��M�cyqH[�
Q�iӺ���^��u�!F@����<�.F��nA�U_�\�Pp��=��O��AF"^w�j��|���O%
�~�� ��궤���¼T,��1���U����%Ǐn��V:���՚�7��k|���L�V��V�����?C2~�����PK5����"  �#  PK  ў,J               86.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G-�E]EG��,��*/���͸yӳ���p���pu��/'G���/;*-a���n{}i������ej>i�x}�߁;듬4M`	t�'�����\�{���*�뺰]�7Llj8~R�vm��'������l۵�Kּ�ȈU��i�c-�38c+q}�U��A���B��sRO~��_�]ξ�gMNx�v	��X�ŀ�4UdݶX�{k�Kg�9K�z�GO$���{���7�q��*��/��c|?�_��������G�y3�_u[�n��<�Ԏ�m�l�w�����{�)F�r��m�W4�/�8i�t�S�Ƣ�xb��s�M���=��q?�x�B��v_A����W����g��Mö�g��կ\�M�G��@W�V�+˶�J>(��SP���+)�������޳���6�!3/4�=��|u���ܝyo���}]tjSS��&<����ե�W�Ůhϴ5���.���.���W/���Uݽ���\�:�d�S^�����?�2'm�	0�';�J(���T�ž��_��,����V-; ��S4���{�2�Wq�e�����VvW�y�h�ɵ�y]+L�45`�f{x�]�c�~�����=u[/U�:�S*�fɭ�}}_�Գ����F�h�m��& PK	�2/  }  PK  ў,J               86.vec�e�a��;���������݅���`��؊���}=2����e>�;Y��\��9�GQ�Q�Y��R�ҥ)CY�Q�
T�R*��U�U�FujP�ZԦNʉ�Y�t}АF4�	Mi�r����%�hM�Ҏ�tHy��^'ݙ.t���AOz�����}�G0�Af���"���`$���2.E���&�Lb2S��4�3#��,7f���a.���(���Y^,�KY�rV��U�fM�b��uz=��&6���l�����Nv��=�e�SA�wP�0G8�1�s��)?N�;��p�s����e�p�k\�7��m�p�{��y��,'��Oy�s^�W��3|k��=��'>���o��{a~�0z����?��PKj.�zs  �  PK  ў,J               87.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG�ì�Ee'y���vF*g���st��z{Wg���q���k���=5��v��R���v�g�s�x����jዮ"<���o�U�r���܂'���<��.l��m�<��|���a�N���_{)�>Z](�q��3g���̙ß�HE�L��Ǹ�GjWTf�ȥ�O^p�����ŉ&]U_���[����KcQ.l���Hy�$��B!��M�=�_�ݛ�Q������%{V�x:[V�sJ�۟�:�_x�5z��ӑOʽVɋ�
�֐��c�7i��!K�&{�k<����

�y/�	SXԥ��3�����j�$Ak:C򅭅z�U���Ƕ��P�*e:+�1A��ַH����&�-����:��X���uG�z���Ϗ���w>X>��*ad�s��#�b���
7�?����%͹۪7^��fP�<;v�G�%a�7�pX�b~����E�9f.��|K��l�-T��ZS���Ǻ87�'�?��IۮLZ��_t��N����B�W��U/5�O��n�`�|�?���=�fu4�~N|�����z�lE>���?�e�E-���u��Y�ڲ�%��Y<����~/����������eˮ(ԆH=��=�:d�b���7PK��&/'  s  PK  ў,J               87.vec҅�Q�3/���������.��.�[l�V��)��dXs��w�LD����;�<�)BQ���D��,Jd)J:��,m��,�(O*����WY�BU�Q�Ԥ�Sn�ɲ�+ף>hH#ӄ�)/��5�[ВV��miG���:ʝ�L�ҍ���gJ�K��܇���?� �wH1T�pF0�Q�fcS�8���&2��La*Ә�
c��Ly���\�1�,LbQ���%,e�Y�JV�:e�Fo����l`#��lG[̭:����`'�����Ϸ��; ��9�Q�q�� NꝒOs����<��%.s��\�:7��-ns����>xȣ,7�Ox�3�󂗼��1���|�#������H��oA|78���_��H� PK
��vu  �  PK  ў,J               88.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG��,,x��q�\;��ڭ���������<6Ku�˘���}�\�9gi�Z��]/�U�GcQ=�=�F�2�Y��Aڵh���{�3m6�l4`�z������mYdV>O�Eos�xqބ}	��̙nG��J�c{ŏ�^����n�E��ʬ}��?+�>�Ͷ��ˣ�&�ui,���ٽWykgM2:l����p����D���+;��l��'A��k��*��O:Ro�� �b��'�Z��g#�t����:���L�����/�s����7�G��3��l+���w	����.oyu<ya�>��WW�X���zS:�C�����ĦU<�8s���~K���@Wf.�E���n���RM��?׃�%Ο��@B�|o�տE����s+��_az����e'/R�6�H 00���W~lS���r��J��?��^nRv��y����;�i��y��x�Jv�p�'�,�.�f=K$�U��|�է�'.˛����k�e����L���n�/��ߴ�:�|�)�kZU�ړdB%��ֽ�*�ֈ#����|��g��/��Ź����Z/�3=,��A�%�������2\K7r����	 PK
?�  _  PK  ў,J               88.vec��Q��ov]�����������l�[�����{=�p����0��D9��\U�<�R̽�(Ȣd���{�)CY�Q�
T�Rʉ�vUtU�Q�Ԥ���r�n�E=]�4��iBS��"�ܮ�nI+Zӆ���=R^t��;Ӆ�t�;=�I����]ݗ~�g �`�x��,b��F2�ьa,�R�x�	z"����2���H�1�n����2��,`!���X�����e,g+Y�j֤,�ڭ����F6��-le��v�v����a/�؟
��A}���(�8�	Nz�Sv���r��\�"����r����&����r��<�!�x�|�|�3�󂗼�5o|÷�w����g��5+�o��{a~�p��_����?��PK���{s  �  PK  ў,J               89.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG��̏�Y,5�~����{��>{mi���^��ud�V#�9�4��nZaXt|����]��\�A_E=��X�Y\��9�������]'&�=�+�w��s��<��{0��s�q��1[}����
Gf�]���qs�A�;��s��kU��~�b��Y ���A�۱���}���,0+��������oI07���9Fd���7���QL�+��á�s�30X�}=x^�wH�ye�_�:6�/����X�ŀ�������g�����'X��?���q���u��wL��]b��[�#̦g���z��)
'2�b���{`u�����3p=M��0a�I�-��G�b�>����a��=�,����/lv	����ە[��oxO(�[2����I?���}{Kgrk�}v���u*<g�߹�O����EW|�����3Wzy�p*���Íu��An_-�͎ߵ��XvG�%s�U)�Ν��SeO��N�*˙ե�`��.<�y�G�	{�<��Z���<�%\�T�Q��R�����n�9`İ�鹭����m����f�}���N��'��>����]�w����C��̾Q��4a�׵�\3ږ<˙�9��ǉ���5��GG7�0��_��h�.7y��r��_Гkş�u��>����g�������~�=eL���le�����o PK��\�T  �  PK  ў,J               89.vec��Q�o6����n]�����[�l�[�O����p����f&"����C.y�S��%��(��(���,�(O*R��)'��UիQ�Ԥ��Cݔ�<��ހ�4�1MhJ3���ha�RoEk�Жv���:�uֻЕnt�=�E�]_��g �`�8oh1L�F2�ьa,�R�x�M�'2��La*ӘΌT3�����fs��|��E�O,�[�/e�Y�JV��5)��v���l`#������f���Nv��=�e�SQ�;��0G8�1�s��6��i�p�s����e�p�k\�7��m�p�{��y���c���<�9/x�+^{�o�[��|������H��oa|�?��?}�_��H� PK�N��n  �  PK  ў,J               90.i��eT�����Cz@���.�AJA�c���������AR�%�c^����~����q�u���}�y��Z@�HԔT� h�  ڿ@- 8��@l, ����G@NH��O@M����������������������0#�����+^!a��l����K�O@EHH%�L�,���^ )�, � ������Xh���h��X�@\<�M$ t4tL,,L�ـy &)���3�wr�`x>�|�w
��SV�!�x�ϩ�i��98�@�"�b��
���UT��� �o��-��ml����^�>?��~����������QPXT\RZV^Q�����������c`p1<23����������������������˫�ۻ�p�0��g��H�q�cbb`�Å���RL,fl29������8������,B��<��(Y���������B�������� �@��<R p��?��&1���Sյ47����m������g�责S�F����C�W��ė^p>�S����W�ü�]�#i�����vƘP!�6r��#���|�Fx}�ө-n~��iU�͈��ە�B���ӏ���^o�GM(Mϑ۾� �Ol}��u#�l�X�ƚ�y�/q����q^#�0�X�?Iê�&��N}��N���a�#`�����u������:�v6�:U�9��k	��gO�Ks�.�zT�E��P�����Ct��,/˷Z�p��+��6��jJ;aA�
z=S	�y���tL�s"p�5�9���@�Rcv>����&6J�F�����N�� ��된A��,����0Q���&���Z�s����0��g�lP��B��p�p� d5IX�V���������M���C��p[�מ�|�C���ܵ�.yqEۛ��M[B����������͇a|W'���Ļķ��߷6IL���e�}jzw��}ظ֖���[��=�y�\b_~�)^*��v�Rl?6���a�$��6�yS��MUf���+���(��D���$#b_�F�O�� C��Щ���/��'��������MI�1��vØ��c�v���Тc��&`�6�6�
Y?�WTe͒�/�w2	��%g�>#w�A�
y��.U�nˤ�zZ���(�r���d㒤]
Bc�W��g��qJ��\͐��м�G��N���Ւ�G���w~o�^�zY�y��X�wEQ�H�rp�b=4�V/�48͝k5tQ��9��3�㤵 3��Ar��d�e���M���E��t{��'����.B3��dcӑ/�hb��<r�iP�	�����
�̆�"	�z*I�OUr݇W����r�����<��?����2"�o!ۭ��j̍Jg�,^)� Eh�H��3������M����㦨R��t����|yZ��tV�g��/�׎��P�������՟���칣��律4W�j�`�"0V,�G��"Bs;����}��L<�1�k�,���^ޤQ�ם�+�SX�p������ή8$_'���r��c�\�����0��TF�j���Cu���2�0s�h-#��#)u�?M���C~��(�F�V��"�u���]����K��P�\ߨ���,:2�`-�v�o��<�f󲜏�^X~�
���1�p�?�:9�D�|]?M �u��J�0�|Bl�y�۴�7���h<r+�|k(�ZVWF׹����mb�K���WUhKas��$�U.��&�r � eQ-X"��7�+�O�7��S�_�2?|'Wk)V�=�w�
�у#-��F������r������g	rC5P�w���t������Q�P��p�h��	��=N<9�a�G/�gw7L'c�M�bj���K����Į�o?9U> T���12My��oq�7Ⱥc�>V�%���!Ĝg{ɝ��ey�-Ҩ:��*g�R4��'��6]����\��A�����cj�),w�mEk��լ�w= �So�T`���l��q�4M�{�L[���^tN�T�*@>�wq�,�`a3#a�ѾI��,��p)���K�:vޔ�Hf����,�m�ė��Z�O�8��P��<SkK��)Hvl|[C}p���K|H�F�O��np��G�H��C�xv�8��J�ۂ��)b;��F� �wYj��q_����_�q�k�_��#�qk��ߟ�+ko��dm�M!"C��`��^$�x� ���R��q�k�����6.�]S5��k~3�BF��݇�k^�_��ͯ��
��gEGo^V1���-�Z��/�;�v���ҙj?�G��P�,Y�hU{D�p�]��5�eɣ�)>�3F,�n{�Bg�&4���l)�8G����1��6�.�	��8�;� ����!������vz*]��2L5˶T��
&ic�o�� ̨�O����<��uh��c��V�>b�!��t���H/��P�>�3ȟ��A)"�����\��r�R������ͯ�0h�ZWJ��FF���U�7��5�J�ǿp%��5���T4j�\ ��Qy�o$���h�h�h�-悡aj�g1a�f(��r���ڃ��Ǜx���j�z���_�W3�<�x�)�+Q�\d��jOJ�_B���*n�R���%��V&��:A;�N*$�L��t^�Boա�Z�y3F��z��u���������#�y�9^�<j�	���E�0n}`�_L49[Q:{<�ந'ݗ���10�+��ޡ ,�Wqv?���-�>������wx���잯z�w�s��g���唴+��t�r�^�$a�s��PP ���N��Y���X!�$�cJ��l��t����c��Y��b����dצJ� �8���g�3pU�ůD�,���]�:sZ�N�l��ʿ��!3y�/��F|���ʮΖ0�?�ޫ>���I�>y��8���O�\��V�
�#G�~��_� �_~+��Z�E'�� ^��4Q˸��?�պ×"�֤]�	�h��#,b�����k��;�X����a�d�X�׮7�U�I-_��S�2׳����w������5��u���I���1��z6�4���f"X5���u"s��fg
�{Cw�:�묻I��@X����|ۂ�(ir��d��}��rLp?4�Q�f"*�����3ȅ�H[��.�̻�*��G-�U۟?7e�dx` z�������j�?R8Xsv�E�2���'��֭��-�o�0ė?�1��R��yi�%8�<�^m�+e&ei�b��~�:�Ma���%:�h�A-f�j�_\�i��1|����yz���7�XS0%A�m@��bQ���Q�Xg��[�AͿ_��0�D�*�8��IXĮ(��'HRc�ޟLT�Ѹ��ԉ�G+�.�v�$Gʝ�*�G�?��#c[[>���˘/�Ԥ�b6֣!
����,�X,Hz�
������/Ԍ31ޛV�N�C�U0�O�ϊ�ĬD�jJ���,�����0\ @�3�����nI�9�0j�RM��)=�qo��Y����fk�<y�l��F2�������؟���+����������h�� �:mǸ3I�J�d�;h�wȧ��O'Q��'��f���bȜ�F�z{���Y-(��,��\ᑩfb�o� g����9�W��4%��aʓ z^S����
��,V��H�D>63n�Xs�N������=���\�
���	a�������;}������)]"��8MF��J�)n��<��X�����|�Kp�|��K��!CLs~��������ML\�U6)1p�<2����U~�݄G��|v!��R���"k^6�{��y1�:S��c�����[e��ΪS�>,z� >L_H��Гm��,2�?�b�$��̵���j�xZ$T�0�p�D�vm0�zg������p�;6���j~�W��Rc������Na�^ݤ����4���V�ь}&�GN�\Iũd��/�ܙV���m��d�2S�
��s| �f��D�/s`*.�~�^^�����a�.^�ӸA��]�D�	��B����rS�"#1����0�AA����Y��D��Ș$t�y9eS?:�5�g'b�� -@5�/erw�Bt<�e���!`�~��\,���_�m��h��Ԁ��!���Y|сX`uDm�}�D`���� ��ۧ{�S
f䈴�'W/�D
�:����gB�^뗞�ȣ�[�_9���]�g�N�,�C���( =��~Zd�D�u*{n�k�E$��lޣ�q��U.�8�/�{&t0�8�K�����64*2��;�i%����"���hwZ���]n�_���X�n���\N�>ƕ~�r?��Nˆ�7:gu�Z���G6�Sχ�9�1>s�z|��D~8
���6�&�t|*��]!��T��i3I� �0��sd�~_S�/�q�/b] p���^oo�5S` .�C�D@�%��j�ŏo/A��OM9E�ү�ջ&�Wi�3���?r���pM�|���A���X��Sp_�2�gPW�]\?チ��4o}�T,��c���g���7�(�QR�UNS����B��� П��E��w�{�(��U0M�9��ʲE��f2Zjٝ~��4֣M����	e#�;�I�X�-n�H�Č;�l��#y�'ؘ��W�W�#@E���j��57	S���Z��Q��|��Qh}!��gb$DU����zb(�<�$�=��o��O��G�������oS�t��Y���2�����gڮ�Y�<� jfX���W&O�+���˲N���s�lA)�꼚c�MG�h۵触�ף��-���w���P����RtaDTz�@��n]M)&�=�3T�F̀/�IH�A�D�\���[_b���T.O�<�]��>�q��Nߓ(x{P�5��0���x;��5�(Pe�>�^T�W��B�,��4�A��F��V\Uʋ:%��_ѷ��j|���ΛV���$�Zl�R~
�8��i�2�3nO�1� 4�Vf��ݏW�w:S_��g����&�s'�[;�XQ�2����ԁ�%! w�鏜1I�-�	���'B�¢���5��L��d�> "�8�@��]B'm�!�#DC��~�슴�)����P�Qw�w���&׭�[�)����E��������ƣGw���,S	d�}�qS���]i��s�����F�d�S��n�_Ԑ3�����p�f�"���0�ؓ�q�d4'��F}2��7��0�\�e�儞op\`���n�&���������G|������Ӂ�1M�d��"�z�#h�p����O��|��p��Su�ҧ��ZI ^��7C�����f9�Y١b����x܋-�A���O)p�Ɛ`e���.���^:�[�:e� p<+RMi3͆S62>�tbo��J��ϔUX�&�����,���iЀ6�O��Y^V�O?%h�� �5ք� �ʾM�Ra���� �uL$��Yg@���C�t欔!�&G�����ٛ3�w�3'HQ�!FX;7墰�^�T�s���XFX��8��~b��b�4��_M����t��u����a �L��d���Q5~~��I6?@�#h����Q�H��}b;�Q���y�`Mؘ}�C�4`��r^�i��<^��`��~1�K�|�)i%q����O�?*�_n�'�\�((C��;.O��s~}�+a���J�4m����y[�}侯���r7~e�R2�;�xQ���C���|�3E쒑�I?} ���ϙ��-ܚ? �Ƽw���7r+ ������
�B�כ!�/� �͚m����J�'@?<��w�(���-_}�uy�V���vOM��xW�J .b�;0
��W�if�10*�yK8˃�o�gf'�x�?(-��A���zgwM����D��J��=%O�p������v:�2�Wo�t_WOx?z#p�d4������Zw"���>)�<�9������qf�cS�)X��Xh�A�UԳ�R]�v8��>��qݑuL=��x�&!�f�S���L�N�>�6�Ł��Q>I� &<:#of�<��C3�����w�8ɺQ���؇���!=�٬����Q {vJ��a`�|���6��� ���i5y!�2MQ�z?�Ls��9�6�[$m�v}��4����؏[� ����^ /������3�� }]ܮ�
",T��:�>���F��߹Ø���D*�!�x�$���(���,�C8&47+����d���.ʲ</ݓ!���818�{f,���"������G�w��14�O�ƂVn�A�uE_C�_I�H��4�T�Ɲ%��(�~] /�X��L�v-Y��vw������4�Փ�zy����XZz��Θ�Y���m�S�0O�x�$�:�RJ�c.IGc��1H`��oH��z�8p8��|C"���o�f��r��F���|��m�no����F}�ł/����˲�p���-��Q�k��E�,�$�ϖ��!{���6�Z!z��:�c)_�|�PgV���l���e횣[۰�9��9uE�K�������S�&G�'.�~�sk��7g���l�����xĩd�x<��9l�,g��.f�*c��G���g��v�2��X��W�y��a9�5�v���]�9Xmݠʼ�� Qy Q�v$��xՒ�sR�O;�*Vc8U-�_��W�q�:%u[&!FZ�>Q 9�ǗcPj�M�g7��'�n:����:�1/�߆9Ҋɽ��_~��$�۶6�|�I")�gūH���4�^[����i[�D,�G�؎Iض�Y83M_��?6��G.t`j�q<p�{t`2����5�4G($�땲�3fz($S����火�H�E�5�}cy�������'����ow"O�ފ���s&h�W;�e]��OVD"E�Q��u�����ڱf��-V?e�8��r�4��^d��&�\Y9�mT�oU���xk!�d��SRs,D�0fD�	6��nn��͗_b0��o�N�	�>h�I��і�����X�N�/�.]+�����"���n�Q�=��(1=Z���`0d����|_'l�:�s~��Tg�C(x�!v,��QI�Md����Xl���ux	�D�;�<�x_ia�:��m���c�/6j^��T�QtgҎ�i|Z&d!Lp�A>���pe4H8Z����5;=1]0.K�*ѥhҿy��|�LH1[�s縨 �������e��J@��~���rFq��jrI�H�yf-Nq䵙�hv?Ü:C�A���	�ø�3A���T�:1P4Lg�zZ���{������9��/@�oq�[5ê�����Gv-u?W���s��L6;��>���j�P����XK�����M�L_��tFz���+�M�/��H�qwY�pQ��ٗ����Gv��A+cm���Ō��[�ߗ�$�
�w������'os�����'E�|��Z�֔��Qp���uɐl@'u�t9�F�����䀎j_�X-�m�hx�T��;R��˹-�I�CN�IK�_�EP%u"
+��7��e"�*�ok�~������ݯʠ��<\��z�[Y�{4��Y_V˟M5tL�N�'U>���I�B�aC��B�+��o�( ��ݢōn�tȞ���ƭ:}��}bkԞ�����O���2҄T	+I,��v��F\7�8*�z�,u�L\�0�Z�$�[w�J,b?����|�0�
�	J�������P�[f����G�K�A�Y�^9�~�e��8[]y�tqXYo�	I�����~9�3�>&_*�LЖ������q۪F$K��//yt [ٴ>�AiO�z��Ƿ�*",�����2"Sw�ۘ���v)s�R��*�����K��
�Z�!HKp�c#�#K�]T�08���pGv�Qüz���"!�<��ReMDNIFas�� -*��.�����zK�n/�4�v|6�J����։ĩ�:Է$&�H��vK�YGq��u�BD�V�"�^����E�XB!V1�[e�\6�ּ�Y�����l��PORa��O���y�0%i>��7f樤d>��1%^�6j��풃>�9@vfx��2��4�8�� �''�|d�n-����ӻ�!���I%����?|�I�N_'��D$�=占�&�#wI�HFC��t"�d����ڻ�qH���Ia ���Mc�|&���̔�K����h�%2ICT\o6�W7/�q�D��.���i��4	S��Lۋ}H���]z|
��n�e�+��͗&��M�Yf��b�4g�b�V-2���|�K;J:ij(}jDʶ9)@��z�e{s'*"2�N�򱛔�_i}|����rT{�bd���pY�ُ�"�:���u��5:�gw3&d�,�E(`�I���[m�Ia�T� �sxP|�F_j$x�%E,�H5�[ݿ���-��Le���``r��}CZ�%uGf��I���ɹ�%4J�hW9߻��/h(-m/����L�jD�e�|�
�-�r:���v?K�C	
��3�Q���W����z-��]�$�/��@+�/a�p/���Jw [9Q	0 ���y�f?q&�[�a}�0��1��������v"F��#
`:g��>��n�,9�N��?�eL4���SCxQ !�O*�q3�F������E��[�/Ѓ�)ytesbs
��e��Ǥ�3��|����W��&إ�m�9�r��?P�m`��t����'Ȅ2Cc����a��1o�k�*<��q����Uy|��S�LP��PK	�"  G#  PK  ў,J               91.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG�(&��歓M�{���?��W�d�O�n�d�7{��ϳ%Qm�s�n�����S��Q3nv��X%�*3�,��Q~�a����?ד�<�e�z����S�">O�x�i��1���9_�ŔN��9��*�ゃ9+,��\�ƾZ����מ	���<c�<�t��gv�+9�7��i�Uui�h,�b��_~͎Xxu��q�)��*��Z�P��6{�5ݥ�>k&��_,|������;�?��˚���[�f��:�òz�Ͽ��lM]���=O�����/*�ڮ�I���z.�`��'a3���"/�J�*a��?�C]��45��V�Et�W�s��T���8"�q�ﳱj�Ӿm�Y�(�{}N}o�t�A�w��������X�aQ��\}�j�S�u�ɵ��Z4����6\���/(��xǛ���U�W�͚v,��IƢ��N��6\^v��GQׯi?�e���8O9��=�ڇ��Vw4�K��XxҾ��Z���w�����)��n�FW��Y��P�Ne�c?���������eož�~l�ʸ�$@�a��S�\�툞��& PK���>�  I  PK  ў,J               91.vec�e�PQ��f������������l�[����8^�<g��ǹ7"����C.�ȣ0E(J��,�g)J�%)Ei�P�r��Bʉ�YD%�2U�J5�S���J�Q���u�G}АF4�Iʋ�z��洠%�hM���y��:��Dg�Еnt�G���K�M�ҏ�` ��1�C�c8#�(F3�yc��8y<��$&3��LK�1=ˍ�Lf1�9�e�Y��0ˋE�b���e,g+Y��X��F^�:ֳ��lb3[�Uo����d���^���دw@>�!s���8'tN��8��r��\�"����r����{�e��w��}�G:��'<��y�K^��;�1���|�#��̗� �Ɵ��7?�G���gJ�K��PKF#��s  �  PK  ў,J               92.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG�(&�ٖ��{ή��f��u�ˉ3T&���\?b0�Cs�����G=��<q��H�@��̸�"��\N^`JN���'���ޖZ*tMh�Rq�xu�_��	��_{1W�u>Z~���������|~Uy�q\����C�g����O:��dq�?`A��uz�s�o����ک���*��%W�9E�v/��Xp�A�����B�����|��H�rƋ�BLQ-�Ƙ��N���&�7辉Yԥ�@ȋ����Z����@�������m\�[z�+��s.���[�>ozr��%�Ş9\Wi,�q�Kc̷��t��+�����=�U|u���mw��e���,��N�����ǲ��N�/������X�D�d��wcO���Zo�����kѤ}��/0�^��α��Sj������Uݎxa��E]�N��W�r�m���SX�H*�3e�rD/��c�6�+�������^`.SǕmT�~��)����CүN��*�ֈ+ɭ��U�|�EěC��Ȟ���n�����w�}*��p��Â0��O+ue'�=� PK �_&�  A  PK  ў,J               92.vec�e�Q��wwww��������C��Cp������9�����tG$I���P�,E)FqJ&Q2I��\�2���@E*�yQ9��"W�թAMjQ�:i&�zo=�>hH#ӄ�4K��\��ܒV��miG{:��Q��ܙ.t���AOz��[��ܗ|�џd��$���Py��HF1�1�M#�%�/O`"����2��i.f$y1S��l�0�y�g�ٷX^�R����d��o��Zy���F6��-l�=���vy;��n���}�O�}�C�G9�qNpR�y�3����E.q�+\�׹�Mn%��m��.�����:O̧<�9/x�+^�ƽޚ�x�>��|�kRߢ ���ŏH��W����şH�PKU�$by  �  PK  ў,J               93.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG�(&��֭�(.��A����uمǴW��5:qʬ���+��vf��ri,��ԥ��	�}}f3K�G g��R��Wc�k]w=x�*��ng�x��q�ewOI��ڋ9}я�߿�7?=3�c�⿍���3R�X����ۯ��%r�<q뜟``?��R��E>X�MYtd�DU��|�a\s�Ym���	[�}�����y�V���w^[�k�ԱJD��|�:����-_�y��]�V$���@��?bS�n�b���9BE��'���\�]'}��៹
ꅁ��w�t��}�Y"R�s�U�H�+>\R�xEq��YF�zJsf=]"����]�Eo/1���qg�%�̟��^��� ���B]A�W��4t4u1��7�������s&��yK
\���U��k�,��b��3�!v�[�y��_[���c�bW��i���jٰ:�_Nr�������N8o{���і?{=���f,<���i��p-,az%�@�)���]m���j���|q&�~��,U�+5D�2T/0=m~�>��G�s�F�5�^XH���?��ǧ������� PKcyp��  9  PK  ў,J               93.vec�e��Q���=awwww뱻����[�l�[����G�K�ž>��a�e���C.y�S���xʢD���.Ei�P�r��SNT�"*�*T�թAMjQ;�F�[Wף>hH#ӄ�)?��5�-hI+Zӆ���}��`�Qw�3]�J7�Ӄ���e�[������?� ���!z(��F2�ь�k7N�g��d�0�i�OL��b���,f3���c>�f��H/f	KY�rV��U~��vk�Zֱ�ld��b��{����`'�����/����;�r���(�8�	���S��g9�y.p�K\�
W��unp3ˉ[����.�������	Oy�s^�W���7η��=��'>�%+��Q�R�����O�K���PK��u�q  �  PK  ў,J               94.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG������L�YX*�gn�Xʮ�0'y���ܵ^�>1Ց�dǻ��ܷ3����س��/��	te�'�Κ��{�`����g�<^[�ui����!�WxJׅ���sk	�q$�ev�Z��|��oK3,� ��_������nۑ�,(��wM�����GK%ʎ��������l�jҙ�.1�]�OX�]=�+�˥�����ؾŅ�t*mE��U0�_�i���J�9?�����4�`��X��M�-��W�ڵL�J�������io��N�����Z"�'���v�+=j!�y�]�kw�S�/�
6yq��.���B|��b3<�N�����ز�ٶ����}Q���'-z��Q����w���4{4u1���?��>_�ɛ������g}?�Z�;m7�ت�oN��r3��l���,n�?��\6�㬭�I���â.<�9:z{Dj���P���=�f��?f�紂��V�k�o-���me�ӏ��]EB��|X�d��5�7��U�H��㚇j^{�L��6���;'b8�(:��P�������/�h�뢬��Uui��
=����Μb8��_��4Íɭ�;i<k�X>�L������P�3��F�;�o PKd�WU#  k  PK  ў,J               94.vec�e�Q�=�������z���n����V��Vl�V��S^9.���p�}f"�,�?y�(B>E)FqJ�,Jf)Jɥ)CY�Q�
T�Rʋ�YD�*ըNjR���I������4�!�hL��,�Gs�rKZњ6����":�u�;Ӆ�t�;=�I/����#���~�g �`���Py��HF1�1�����xy��d�0�iLObF����,f3���c>X��(ˏ������`%�X���\�:ֳ��lb3[|��v�&og;��n���}�0�;�|�C�G9�qN�4Oq�3����E.q�+\�׹�Mwp˼��r��<�!���c�	Oy�s^�W����-�x�>��|����(�o)��H����S�%���PKs�r�r  �  PK  ў,J               95.i��eX�����YT�a���[�A:�CBZX�\�S��X��niXby��ύ/�ý�̧9�<3�{f������TMIU	�� �=��"@��������������OHADH@@HM�����%=�KZZF����<@ZZN^>AAAv1)Q~�����Y��������������Y�d�h2�4f :�c/���Xh�-��!h��X�8�x�Oͤ t4tL,,L�'k��I�E��'��l���A��R����M�=~�"`������KV6vN.A!aQ1qyE%eU5]=}C#ck[;{G'/o_?����Ȩ�ظ�Դ�̬��9ߋ�KJ�ʡ�M�-�m�zz��`�C�S�3�s��76��wv��O��/.��o����B`��O�?r�=q�cbb`�����?d�XL|��`K�g��a�r)�����'�V����Y�����������������Z b�=] 8J��ü�;���&�r�K����J��������㋧�d���*ZM��57�!C�Js�z���WA!�*����՚ڙ��F�N}?�G.k���~�������ܑ�6�K�q�Ph����O��ɏW=�j��'<15b�3��aF�>c�2 �3��s��È������
����k�gf��}z�7�(E�wY�ć���w�i��D�XE�C�[�$���B��`�$�e��u�x�bcG�\�C9,���bY�w�=�5��Y�7��gM�
�6�s�~���� �2�?׊3S���J}H�qK��ث�c�-��u�e���TL2�6m���`�.WJ������,��6��*.9�����s����G��Ֆ(e��^U'�%�ǎ#�������EX�$������H��u��b>�&�X��NBw<��9�<��+8�r?��ӷ���~A�$�������vvJ�C?�$��=�"]�ő�Ћ��L粤�ӑ�!R�*�*�Ǳ*�D��0��i�Nfh��iʱ<�ώp��M���,�m��������et�
��T�I�E��9@��p��5%"��G@`O�©؊��6\�{�ۅ�?����������צ�]2�y®���L ��#�d��d�%
޵�>�n_y���raq7ˣc�T+V��0�pF�n0ɝ�kJ�����8t߈ܠۛ99
�}@��2��l� /��v��T!�^�,�Cf.��~��g0g�C��+��Z}�b����Op�gv�E�/�C`�Ӫ�d��x�l�AyU�9��|8��fn,�-'T���*�ԱV*k\��XS�ܱ��\Kn��8r�5��@�D�ۑm�ܨx������\��%`��`,#�=�ḂbA_��lw�EK>�7_H�a!�*"BCJ]g��ֻݏ ��K���<�%�uBe߳T�W�����=��Ƈ�u��>����K
.�-N<i���?M�zz8|��e�!�¶�7P�[��� a �kK������ve:��X�߯�z�M��@Y^L���iߺR��M��L	��Vl��C-R7e�ʶ2����8:&��%��z�Dىd%r�� � ���?�����r��7(���$s��@cq����@�u�A-m?�B����V�Ol�.�ۃ��3��<:'65�\G��la�H��N���u�Q�&iNMR��O���Һ�iBK��D�:� �w��l��m��҇jh�2pM��0�Ȍ�	�������.�q��K�w��&q9�Fs;�x����g�,�����ŝ�U�L�xTKA�Ʈ�=;��ౄߞn9���*��X»j���u&��t��9}]NB��O���-��Tr�n4k\Am��B
e�mY����Fn�s8{��#6j��@�3]1L/�9�\g���i@�8��e�ǩ�0���ۼ�F?=��_��A{�V/�_���~������@���������/r�i��۬����q�7��v��pU(+����鈧j���k/D\Rb9���>�{����%�JC��o���n���wڿ�5U=o����������,�ʦt4"�ܠ��B�{��}$�Il�)�
��@����g�UIU�}�gO]�zD[mL6]��oളe�Z��DCT�q�I��X�n�$l��]zƜ@*z��w\�?�K�b3��#v�(;���+�-���p
���$�7���K/G�<T��ä�������m"j��p4���v&�W�K�H�|0�1+N���Y�3e�-t���;��˪�_��4����S���nE���31�K?�٠���V11��΃~����s�5 ~�d0֙/��N�i�>�>���I�:�tXx�tט`oŮ��3$���'6�.�뾐�8���8�X�~9
"�7G<��w��f}��LO�:]�$��>l�u�Y>��Eʹd����Ǡ���t&���,��ӣ���Wŗ�=W�%��i��# �.����M�r��{eej�68�A���'�0���W�D�]Dɲ��ͪ	&����Je��Nm�t���K+"��Q�%J#������38JԄ!�|�*������eoO@���űDGŊ�tln�
��s1��6d&ّ3���S��|  �S���<��{�n���ٌ�|��ؽ��K���s�>x��K�����=U�8D���u~po�<e+?x���yF��~l�����,n�_.Nl���9�zr��� t�܈�C(|bL�E���a�*�,���-g������+o-��qA;'U�NŹF�mwڛdYR��_^�\��}�Y�_��J�,��V{�S�z9����V���Uou�\ �vYJ�L��{_^�9�CҢ��2��[�b��v�6C6�t�rx�LU01˗g`i2��] pΧ������s��D5姅��_?�Bնy~�X�TMk�8���V�w�CH�t��+![M,�
7�R�:5�n�StDN�c��т!Tӂ�-9P@�HJ��ܔH[H��g�0�Ϩ%n۬���Ǚ�[$�>l�@E�.�e���H\�[��S"��<4kǰ��X��a�r�u 6���<Y�vW��o�.���/pn�]���S��X+��By�摏 5��Ҫ� ��O�� ]<pR���Ş�k��ŧHۡ�MI������V����ô�0NP����4�xFi�Ֆ�"k��KG�L�4�$�B��b�O�æ�?��Pm�z��=�����`��S^���l	�d󇵿?26T�~0�26u4��S����D_lP����t~���z��B'E��,kv���T��sZCT��!N+�4�Τ6��}l�t��m�����X*�_�o�sQ�Ξ��� ��3�>ܳ��"��S1P�v�3����EV��T��3�.kCw�Ś�Р���߾�_@�af�q�Fof��┨,����>�z�l��	Q����.���=7aV�����~�^��.�D�;xA�k�����)%�m//Z��0��;�sO�珀�f���R�Մ{̴�u�7���5ջ^�D{���&FE$ǏASpX��<5��;�ޕ=x���ޔz�4�_���%��:�OOi�������R3�؍W�_�X�@7}����58�a��v7&J ����
��P��L���,~K?��Y�^�qW�EQe�� �<��s�~�2�L�l4���=�.<߁Rj }�!�,�pp��������T]�E޶�y��5�V���,1�;f|L]�i�5ueC'��![&(�!�s-`��YD�5���r��(������a���gFe�M����Ku:ڏU'�duZ�H��><_��V�Ax�Ig��j�kd����	�� lg�A}p�[:<�CL����Z�|��S��|U01�蒊J�rS{�:Ci�W,崒�� Dd�����/Wy�$�u�g���k>���̊���Nt�y�M����f
���[p�ߖ~�v|E�Jm
���;�����e���x�*�ɒ���M%yU#CNB�1�o��Y��.��iq�4��O��V��:}و���0� ���1(w:l����z6��A�؈?���pw�,���,�>�ҭ�}�V��.͟�z׆��Z�	�V
]*\Z �^��x�n��׋4�M�}Ϫʸ��c��!���Wj�P_{CI�2A%v���3���.F�B�O�NE��%G�?�j%����+t%]���9r��w����ҾOi�7��� ��R�4e��K�O�|�*�+䡩�93cq;�lG)���id���U���?���� /ѿ���m�Hz�C ���W��|�HAED�؃JUP��g�b��D�����*l?�O�ӏ����e�o���1}�S+Sc;���j^������i���l��yw���s+I�/�2b�����c\��B�ݖ	�ޅ���7��uu������=�e����sz��F%f���)��F�ҭ�눹 q|�C�Ԉ���$Wb���X��Џ:���}N���I"�CoH�S��"yî=�G�+!WQ�w�ulc�L�D�����Qb�.z?�%|�C���A)"��O�
2o+��	�ZF3�J#Ts�)1��ɔ��iPq�}4��@d;�������@�	c�Q����,�/�c��� ��͈�Z.�A���B�2�ʲ(�xv�M���}������u#���H��69I=��QqI�	L�0���6�r�ۥctY�Br�9x�rȬ~W��2�f��@f�4D�l�]A��E�Y<C��{=\n�Ko �h�(j��W��h{��ő�Y��j�02��� Q�U�־���Z��$h���;�W��l� ��j�6�p���;mCզ'<��h+���-��aԠ�3�B����[gGzQ���LEG�l����j�G��E'}�yB��	�Pr��y�/��^�¢��-�W/xSw�u�}��&]B�ȝ A�p`L�d���t�Tы�	i#ʌ~D���+�C5��n�^��SP��}X�B�}��s���2�6d���oY7L�ogD�
ˆX��[狖�Imn��<?Wk�R��
��l���_��6,���=;�~YI����+?�B5+A	
��hPdГnΔ�SƧ,����]����w�y��AK���Z����2j�L�?��UX����dTJ�  :c� ���/]����EBlU�ZCExl��.;�S��&[	����H����y�sA-����c��:*��i�S'M��N���9��N8��/���Jz���q�	$�ThW�~�KQFm9J"�$u���%"�pچ�H*���5Y����Tᗧ2�� �Jc�7����C�\0��Z���nD� ����T�<�(�V�a{*���JzWw[�}��VY��G��tb�0��>qr����kj���*����*�s�\��j��I��{��cdd�.o��b�2�7knnE�9[�$� ��ty�#�¼����CʹEHW�µb���d��W�*s��T��-��B��K��^h��=�lo�Q���7.� D���D��T��a�����e{l�uRC�J�x��,�ըۉ�&�܉�����(��t�B��\J�Vw',�AF�n�d���>f�����	(\^S�jj�pK�HL��$0"�]{p6y되17���d��� �|ψ�hW'Y����Z7�(g���<9i��[�$菠Q�_�r�^vnn�Vq�J�ե��2�����?8
�{���#�|����X�$o��D	��&�2Dz��5!ב�+���};��.�jԑ7o�/\V�((_������|��A��pq�Y��x��/ތ$�=��c�H��fF�*�[b0"CL�S`�
h���K�}aq�����C�A�0=u$1�@ʿVj�w&,�֦��k�z���� �L���~HHq �m_�d�s���zj��"!G��I�4O�"�6"��H�6{��K��������l� �$Z1�|WZ#��հ�ٰѪ�g�3��h�Ñ�M3��,��P˰�F�� k*Í/�	�&�C��>/���Vt��d���(��75���V�[�J��R�*ի	i�X�x�� v0�)�����<��[���쌥��9�B50�A�Q�۠�#}�`REJYi��l��em�G����D$�?KFP��+x} g�qj��*���,��cD�ծ��T;iK/��t��B�Gn����~�^8�C&�"{��93��3ђp���5�����"�xU9��v��L�	��;:�6�Vf��D]�_�%0F9�Z��qya�?�2a���~a2���1�$�NN�l��E��,�(t�v^3����������	$d�ɻL�!8$z���5: ����%,Y�{�_���or�c���G��ڀJ�">�?�V���nZ�Z�Xia?W�{��@J����Z4�ը8�h�����j/q�SPn�A0^��ۜY�l��7GOau���3������UP�-��<�z���,-Q�x{�9Y �b���u��y��Ap|�Ԇ��a	90�,"���Զ����n~�����<L����|���&!Iy�ŧ[���s)�hU�\v�n���V=xə7�b`_N�^�uw�Q#q�wG<h���_����G)j�ֽ��7��xX�E�}��ڍ��Y8�C���-������$�]�~K�k	{>s-1T#����,����c�Z��j}����t)�Ja��>����7So�3�}j@-��5[�"�p�~>��l�����n��.�gU�^3`�J����ϵ��Ά�v�� �_��M��/E��v%&���LA�p.��e�\�xT�E:�E͓V���_�n���b�a����E9��[�>�nGJ8v�'�'58O�%���~段����3���Q��"���BJ�03��A��+����bs=U�셜�hܼ�?�}��b[�C��!�D����Y�
y;�Z�(:mC�Hc�%x�c,��{��? ?�@ȟbϳ%���Pi�"qLiw���	�5ܕ��W���
�5�=�0M����9���Bz��j��a�X���t��;@7ђW� (C��ֶCqd,>��_�Yp�;��ԋ��4(�ѵ`��!A,ՆJo�Т��`dx'��{+�WÚ�O�*`A�-Vl���e��Ĺ��$�	�3���'½�ı�,�pG*�s�Bu���r�J閕|1ʑ'���E��KA ����p3��(��WkufkV�^,NF\���B�NH��0�&�-�Pzr���Ȥ��
,UƸ�pLD;�ﲢ���������G	'27b�cղn����R����~��g�N��]���J4+M�0a�גZ������.(7�Om�
85+����c��uCÊ#W�v��rA�#�V��d�T��(��][`��f[�F^��/?]�(�	h��FX���7��^��N��u��"!%�����nOY����F����?�ܨ��t3	�-��.�I��~\H)����K9mM��خ����u��qƈ®+���ͮ��aݺ�~����!W�)�d�e�p��P�*'tW���&��w��l��5[r��O���?��E�	#7�^�I��F~��w�Kߚ|/�v�coh�MW��%c�%�)�
T٬��ڕ���r�,�Wb�6��Ak�]Ƴ|K�
�0r�F:��e�-�p;��ϛ��
�%&�,7��O{���_��l� �'U����s�o,��S[�CJ��B���W^3E����Xh�Wban+n��g�{�!��+.�x�H�R #3�.G���ࡥzڤҶO/3�X�W!1�d.h^�؆/Ξi��ҥh�-���V���ˈ=i�=��Jr xi�䥁m��Vq����wE[����'�v�ח�~��8�K�;A���n�5���sW��"�@�����AR��J���H4��3�/xM]=�'t[q-�3����B1�;sZ���j�Sq�J=�I���%����<�*��h�UJ�YޡyИ�IA ؑ�P+�n?(�&)�	�:���OR��q߮?K�s)O��=�ל�c��Y��i�����5+��	2�ذ7�I�	!>�U�_^�ܥz��)��Iw��Y�[���*�������t���.4��}{%�=gA����c,~�x	�� F�7)�A�0G��^�v��4��#=���7�dK�]��]A�(]�q��9t��P�Uƶ�;��[©_��,Y�ﭐĪ�$���N	�iA�[0�8]B���5�9�0E��A���3�Z��KPki�.G�J٥����`�����;6i�ZƖ�z�h�򀛟~�I�ߍEiS�t�ö���v��ia��&����7���^�vr����Ld�E�����w�"b�"�%>hĉ���a��
��Q�)"s3�i�ˈ�I3^]T��
��h4�bVȗ��;v�\x��/�H�q���?�4α�k�lB�X4����kxe�E�-Sc���vV�v�3��H�W������I;a���ԓ�|7�tH"$~��l<!5NKk��j�ݧ~!ahQF����i����.��2��aD�S���KVf�������yOw���q ��h =�u/)�M"C��-T.1��
�_<�XP�򚺛f̦StpV[�ɦ�_�0j"� yJ,�G�� ���K�5��^��A]�+#9c��+zԥ��*P��a\��� �mzX�8ƴ�K�ֺ,�cѶ�Mc������uԳ:�
G�!d\�s�Շn&�` ����"��k٘3��K�HV�s��Q�|�[��o��s$�G �(M��~�7j�}����
c(��*�k����xU� Y�c�#Ì/������6�I�Bj~����#Ӄ5�nR�]���x�e�gh��O�9uE���PKYWE �"  �#  PK  ў,J               96.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG��,]&9_���5DzU�.u�WeM�쓣N����Pw<#��2o7O���7��yvT��E]���"tČ�W2�~{\�A����ua�n�88�ɻ��_�����)�Ȭ���[��Zr~�c���Ezf�l9E_��:�:z�=\(7!$�R���Y��y��{-y�X֥�$ �����1/�t<�a����G���G��Z�0kK�'�%[v���H{�e�^\�-�l�;]O�L�r(�%�hq܅���un��Oʾ-�>��j�MB��YϞ�4~ݳϨ��ʶ�&ui����قw����t���dŁs���?�3r��[u��ᬞK�s&�O9W�i�����]c����C��5u%si,j���r�^��\�p�;qo�o�)c��ű�;�>����8���ꎿ�}�n���Ǫ�r�u�Q�@���4�`����g�m��s��.�<(n���m��|���,��_�t��ɽ!Z�7�����;�̕��*3����S�&. �,v>R��)yh��v���<�}�u��F^�{9�9vLO�1�_ڹ����!��΂ʨM�[槭:�|�7��;K�â��$�GJ�:��G��пī���]4�Q���hp ׬����N�<�S�*���/uMv������+��y�V���=G�[(Z��DN��:�,cQ��}�5L��-�u��]��� PK��N�c  �  PK  ў,J               96.vec�e�Q�=�������������]`�؊�؊��p\2,���a��DdY�
(F!9�S���JQ:KQF.K9�S��T�2U��f���Ԡ&��M�R/F}�m 7��iBS�ќ)-�ZɭiC[�ўt�SJ�Y��ܕnt�=�Eo���W��ܟd��P����Y.F�#�h�0�q�g��D�;I���2���`&�R>f�7G��<泀�,b1KRK����Y�JV��5�e��zs��f���ml�k��Ny���^���t�Cz��#��9�INq�3����E.q�+\�׹�Mnq;+�;�]�q�<��y���|�s^�W��o��w�{>�O|�_����(��?#�/w��;�'��7�?PK�T��m  �  PK  ў,J               97.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG��,Z2�'�^=!�-5�ʞ.6O�M��ܾ3�����Q�G���v��	;��{��<Ϸ矚�x�۩U$Ї�Kc=1�\g���������2��Ψ��E��T&3��~}�G�JE��KΛ?����7&F���6�Z����c����:m�4������U��ɿ��5?��z6+�U<cQ�Ƣ\�*�Waە����Љ��1�
z�w?�]ivƂ��,j�8��u�/�G����צ8ￖ&,1[�L ��9��M=r�<�J����r�)|v1��c������@�m0��Ӻ4V��0����^�%���d=g_d��A��19-3��7]c}�j�&O�S�)��<�u]�3sF��g���Xԕ��g`��f�T�2�H����0����LOj�}��.{�Gg��ȹZE�����M�Ɩ��T����*�E3	$2��9b��N����x������'o�~�ٺ�#���=u]@�ii`�m�ua���a���WWp֝ݮ"A&��mn�t�SM�়}�:�}]�~�m���DS3������˵����؞�+Y~�_���e���(�,��![+����>�Sf��p�=o�Ն�ɧ��\u�$�$�n�^y�i�ƟGV(ˤ<������E]�ui0`�L@����>��΃\�2�qޜ<��q�z���#��|�wE��-�u��]��� PK��[k  �  PK  ў,J               97.vec�e��A��vwww����ݭ��]`�؊�؊��]/.����0�e���Q�|
(N	JR*�E�,E�,�(O*R��Tѫj_5�:5�I-jS���K�Q_��ܐF4�	MiFsZ��h��JnM�Ҏ�t�#�R��z]�t�;=�I/z�Ǿ�z���2��b0C�"�e1\�HF1�1�e��&�7Q��d�0�iLg3S.f�7[��\�1�,d�SK����X�
V��լa��:s=��&6���lKc��y'�������p��z����(�8�	Nr�Ӝ�,�8�.r��\�*׸�nr�;�6�p�{��y�c�'�S�����y���|�{>�O|�_���E�=��G������G~G.�D�PKSV6�l  �  PK  ў,J               98.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG�����M�0G���M��w(���Z�.�~Ym���i�>v�T|[���{�=�;-�N��_i�x}�ׁ;듴4�`	t�'�6?~&�'!��+���_ۙ[q��φ��v����'�7�%�Mp�/�*V�9��0xc�c���ӚY=�Viq*wn�sz����z�����<��9ab^�Ƃ��4p`�W��]�|��N��i�lw��+�~m���G�I�}��^v��g_���x�~̥���f�L�"(�}����_����o*�j�z��ɗ�m�lí<w�}�L���H`�>W�����b���5]���O�G=8&<�͛ts�U)�B�m�������2�9k\Oi,jl%��b;m��<�AH�܃~�g=�Rs�|��G�'�d��nZgd���:�c���7���2�KcY@���x�b�9��"
a!έ/��,�x[����Ջ>�|�/T�%��z������Փ_0�Y�����_�&. d����»g����E���{�Q/���n[q�A�l!���W�͚vD��bW��i�V���k�m\Xt��m@��˭kn�D���x���[��v��0G�in�A'-��_�J����͙�۞/�Xe��yŢ��8���{G��X��ņ;Dl70��} ��9V���OH���k��dE��-�u��]��� PKT��)g  �  PK  ў,J               98.vec�e��A����kwwwwwwwwcww�-�b+�b+b��]/.�����DdY�?y�S@�b�%S^��R���P�r���D�U�*W�:5�I-jS��� ��՗АF4�	MiF�z-�V��miG{:�1���Y�BW�ѝ�����E���џd���1,��py#�h�0�q�w��2Q��d�0�iLg3Sa̲o�<���c>X�"�,��-�����d�Y�Z�u�z6��Mlf[ٖ��v��Nv��=�e�9����!�0G8�1�s����4g8�9�s��\�2W��5�s����
�y����>x�#��'�S�����y���|�{>�O|�_���E�0ŏH���2Ga���PKu��n  �  PK  ў,J               99.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG�����
���=n���������v��Ko�����c��i]��{��4��_��r��ީ��?����;&�������D]�s��g�n��S��������2[�'�%��J��W��}�u�����v�����d�'6s����2T�w3}1OM���e*�&�B��Xo?��_���&'<�C% �U�f��5���$#�S�3�Ȥ������0�Ǻ6{�|�顕�3'li�q.��_Ҏ���\*�ɺ���%O%�Z��BOx��c_�i�^�J�����o���<<��L���H`�¢.�y͵?��	NX�r��k��;u_>��n�n�9����7%t�5��{ll��6�:��"���40��|���7�j�eNs*73�?���:_7�c�M��h�^�|��b�E�k��'�nc�m��1�����RY���ò��#�/bԖI.����x솛B�,M��sW)�!��skQ�Jv�pce�"�˟�m3��L]n��/ۺ��2���O���7���b����v���L�ÂU���Y�z�b+s���e]$���hZ|����>ǯGK�j7��e:''2��'ڼ���-%�h��9���EKN�If\N4N2�&��4�
\���J:-�r�|�(�~��׆���x�-��j�3�nV3��-SrR���o����|q9�=%q�U[�U}�{�����e��a�ſЋ?�^��^��i�9�����C/t��� PK\	���  �  PK  ў,J               99.vec�Ŏa��S�}qwwwwh������%8	Np�a��?�TV�7ةIUD���'�|
�Q�┠dʋRY�Һe)Gy*P�JTN�Q����jT�5�Em�P7D=���iDc�Дf4O�ha�R��5mhK;�Ӂ�)E'�κ]�FwzГ^���>YD_ݏB�3��b0CR��,/���`$���2.���Y.&�Lb2S��4�3#���v��l�0�y�gY��Xl�D/e�Y�JV��56k�u�g��f��5��mv��v����a/�؟���A}���(�8�	Nr�Ӝ�,�8�.r��\�*׸�nf�q˽��r��<�!�|�������%�x�q���|�#��̗(����"�w���'�"�PKFo�l  �  PK  ў,J               100.i��UT����_�!h� �;$� a����]�'@ ���=�C��.�w	&0|���r��[}Yu��������ŧ�����,�� H�x�H����h�XX�ظ$x�88�D�$Ԕ jJ**ZFnZzN**V!6�7<��� �`^1n>~��l�������K��G�KGE���lO� !&����D "�"=���s�!���Ð�QP��10��q�_ �H((Ȩ(hh�����g?�J�FD�#�N�a�A�N��X�� U�C�9}��g���M�����������_@P,,"�NFVN^AQK[GWO������������냷������Ȩ��1I�)�i��Y�E�%�e���?��[Z�z����������7��wv���..��o������Å� �O�?r>s!����b��	��?��ht<�D��������$R�u=X|����d���L�A�o��;���/������\���C! ��Q�Z��^���{8�#�3=�R�v�OS����	 �VPZN���.�PeXv��NN�~���`� ����ꃷ,�T���1����$[�Y�
��>�ר�r�z[�K�4�s�6�jȳ��Ty�"��	N~?<�P,T�Ī�	xO����[xU3�ǰ!H���<C����?����ۣ��͇�"�B�(D��`Dj�V�"��ɲ4f�~�}�*��T�J����M�[��P/�a�.u��q��υآ�\�J���yAE���Ϋv�F���?Zń��^~��H:��m��q��f��hy{<ů4빡@���H'��6�B�g�;{ۀ�P�
�#d4�A|C��� n��{RJY���*E�׊�$�#���J)��-p"�q���F-1My����F��XmR��/�9T�h2���i�Y��/���ĝ� c��'H�|W��������J����ԛI�UmwL�C�;��r����bZ�|��ȣ?1������%X%�������;����/��//�	D3���Ht�P��|[��,z��~�?%ߐ��2�
�W͎į=�6�Ma%���6���~�^N���+�T���J}���K��|������D#�C��2�
��E��2��5Eu�>m���S#M~��~d�rF�~�,�6>�CG��1&���U������UN��v�!�ڟ1ϟZ�����ӿ� ���hE�,Կ�����t	�
�4h����>�L�*��H�{�4[(Y��`�_�V��/J��%�K]�8فi����_�.�ϗ�}�����2���԰�gl�=/?��a;�C�Oa�◖����y��>.����?�'16k�D��T&.���O�]��aT\�����@��),�#r1��p��
c���-O�د�ج���o���{�����(e��/��	�U��O
���C���ё�-�g�y4V��my4ҩ<�^\WX��@?��	�h�+��"1���2�(lLTǵ^u���<H5�Lu3Q�7dVZ�����Z�����|Gl���弿��Y+m͚�z/�W�*h���V��s�����r�\T�ev+��8�k��xb:=Җ����?¨e,�A�~i�͉{��Lݳr�NZ���l�J����Ҵ���~��$��n�i�xGop���6��CZ:ab
A�x��l�ß�5*�t�so=�����Y
�h)Ǉb����^�4 ~��c�I��۩�HM�u>��h��𭨩����gC0j*0j(�@�,��y�����MW����c��<\�;��5%�cK��
%�[W��t7Ї8��|
R�V��U��|N�v�W��"�C|?L�c^49D|	(�Î�.�g�' G
}�tT�[Z�_����z��a�MQ́k��ko�����ԺA��M�4����?����w�XL��B=�����+ܿ�1D�#���i o_�F����*BC
���j|���Ld?u��n�Y���o~��:iK��7if�!7��UY�s 1]���_���g��N���s�bԓ,�rh�h����'�)�1���b��#�6�!�U���7��.����x! ��?]�p�q|�lݲϵ��8������ޤ)�&��*F~��S3�2�8:�2�q%.nCH-�0Q.oQ�O��������?�T�j�Z�F�S~;[^r���`Ƿb��Tݞ��Hy8T��I�0�Q�(��)҄Sۇ�*L$�Ykd��Pŕ�<�xp�p"��Hb4Xq�QSHߙK������r2�h~��4e�ANF�� ��́s�b��`¬�R����G��� �������fM������ye�̿d�|^���L�-�-��CinWHY����_6��n��#2�u�#�T�v�ah]�_z�4��&�G_�F�-�÷�������ڱb��z��dPJH�v2���c,���O��<��������_���3J�v�i* ,lr,��%V�]�%{�+ꂅ� Ex��<���^�`����0��dyCh���)��
 ��K����E�('�?��"
B`�0v,����K�h�a�1�i7|���{��T����z�!�ӓ����l2��}z�i8�y�֒�u�{�J&؞b[ª�����v%�l�&4)����5�u����on]��2�< �L�S��2�*O���>Tmshf�OOCx�K�_��#dj���?�tK�	i�n|L��mM�*��A�(4�]%L@�+�����d=�n�����zVdi΢(1KFL�C���-$Q��*sW��A�3�`�5Ft��X3V���ZO �����k!GN��"B�n��Y����(�B���S��5� -{��ۥd��z^��!!(k�^?��]���`j�H��}��PV�ג�&k&uE��[�wp$�T����&'����$^Y�r�A�W��������>
�1;J��y6�|M�kx�̼���4�S�{�&�Ƴ���*�a���ku���4�����U_�Z`g|	�ϴʹ�3���B�LF-
�q��z�)0L�T�Ճ��څ[]?QQ&m���oʫ��;1`I鰤�F�[��#}����1����eM��l�쀾<ŔĿJ�I(�9F"�_�Ɠ=&P�N�PP�V;4�7��kL�ʕ�)+׎�,ȕ�;��`1�"��V/�m���^�;jF��W;���9`�KNny�k��ԷB��\J^�%b{Nz��AR5l����uX�z��ٙr%��a���'t�׌��4����7�D}��{FΙNL���[nL���������?}P�0��MhYY�[�p�s`�S�w�P��31���={�Z�r����^v���$/&Q��i�S��DO־�W�Ҁ��K�H*�I�kH���ja�Z݅<�%9%��l���3�佮���kC�$U�����t���3�C��*�:;�8�/8�\���%��х��=�*!����׆��|%�+7|�Y8�=!��·ƨ���1������U�Ɲf�Ã�ձaYM4G�"����fТ��Th�J�IO%}��	��K�{	���+ֲ�ԝ���Hf�L,��f����&���Ds��m��v�9�e�'�������"���O��M��V��q-������ł/�<nҤ���xiȼ����E����B���/������v�L+<~+��'��	X_�Zi˻Zj��,b ��ZI�>��em��K�Q̣�A��>4X"Cӄ;�cu��&��Ww�!��ڍ�H���t��r�c��G�%Kl�}��C�\�U�v�:�Ũ.~X|�~u{r�}��Dϼ�S�؜L�"y�rlQ�zt�X/��F�7��^��91B�����"�	�t�.1��h�¦{^�z�f9�����	��03K�U�E����9� Et�=	�	u�' t^qD���P�����ä���V�ွ�T���!zh�)����3��z�5NSb�w�\T�r��
|�2?nr�,����t͔:�佻��].���ԢH2�O+�ȕ(.��޸�$��{�A5%�����&L:;�N�}m���6-�6�!�	�T 5ަC~�I���h�[m*$x���K�o�
�nnz�#�i�{ð ���(;>�L���gdj,l��Cc�^�׼��
���`Doc��
�K)Q��$��� �^4������9v�~�UMmx|\��m�����!mYϚ�O��V;}vu��3�����פ�+2R�l3�FJ�H����$���@�,O�M�w�S�h�0�ͽ��ʰ���8�����&w�䑣�Bb~}�nn��f�O������_��3qՉ�����=��4�^�IL (]�F�����ߋ�ء:�w�O�`������D�s�~� tó�	�#Y�<D�*�C�^K��\���ߩ~LLTа��˿Ε~M���3�,�,���%F�U�F?)#MQ��Դ��Oܒ��/��c�[�z�(s{�����Y ��#�!�93R�0�������F�^��y'�7<ka�H��ė,n��8�r���(D����$�W�;lӏ*%��*�t�]�~���%�"Nk�(;�7�O]�Q�xDp�W[ۇ�?�7���V�n��/P�E����=�zr�:̨���$g��uU����d`a�ʃ�*�K���}3�&
Kj���4�v�5	�^j������>�]�ߛ"�/^rrc�	h�n���u� ڕ��Ğ_?eQ�"}'��FA:"ŋ.�E�z�Kl�`�T�eb�w�o'w�e6�[�m�		�a�h�x`����_�V��������?��њT+g�7Hx���/0����-������/K�^��#F�r<.�C?� ���s�V���:����g�qQ}�.MV��b,��+b�86_�71��O�Z�\D�7�� #�1�Kb��6!D
��o�����I �����!e���j�TH�}��\�d���d�2'�忬��s�=֖u����a�#��q�|�c�LgN\�Р��t�u�������gA!�d��}��,`��ۯ�ț��L~f��D�����9�����K3�S�:�i?fe��ㄩ�#�2��}���L���Tߊ�9���!��n�7 ��p��$y�eu�n�F�޾~dgi)jMF���U=�������\�ѫc�+�y6���m���ս���{�rޙg$�Ix�p���w# ����b y���:X�J3᫤�������;A�g�]pXi���Kyb��t,�{�΋\c��7Nj�rzH�VDS'��?���ʦ��JS�8ߐWf��/���;>�K$M�@�����p��s�:�o�8�S����s!k��r�b�w�'�N<�&S���C��U+�Fb�)&�=�	�\�=m���*p�tdB�k���},[anD�e��'2`|}%��P�4,5�M��s����|�����$W6n`(37�_F�GaN7|k�P"&�pgh�� �D��T;2zM�����oa�J-�,��.�r.9�_�S����"��o4�f��0���%���
�0�{�z���p� �'��]���M�H��g��O�J(�6�r�؛��8�5bF�L_$I�1��`,fnv8P���Q��'�7|;�0g�
W�|��������H��bf�}����O�QJw_4�%��0�꺆Z�=�iN�ݗ�
��.��)�Г�q�OR!�=�5��s��벱G�?w�u��-�"˿��X��~����N�~l(�foc�h�|�)�1Yy��r�h�:�,��J����*u�mφ"�����!S�8�̪w�1�C��BU��ڋ���Оr��/�j|Ul��:J"Th��)�Gޥf�3�VkYr
Q$c_�=���(���PQ��x��e�V0�6=`/*���`A���WX�~i����J�\���5�u0����~ֲ�����7�0G�o��k��9����ޒ�}E\��:SwR�U ��s�~P@x!�S3K�
��7����Zw���T�t������r9K������I;|	��e���1˟�^���T�K�h�^���ZK�����2W���tuJN땲����I6I��N�S�HX�܌}$��b/�4&jyr�K��d�0����c�:�.hT~5���Z�HM��uυ(�.ZB�)���ŭ{�qZ�Y���K,#�`�!B����5;}��|�!��p��詧�*�Л�ufe	�����h��'*���l�B�d'��'??�۝��wJ?Gvh�t|L�|�J���ѐ!�>x�4���N80�	�\Ll\H�C��˟��7g�ӡ8�m�-g�Ar%��<�׻�������$�k�
�f�r��i�8�v4 o���(��V$!v��as8�-�����?���8��P�]ll���{o6��W��zJ���r;o��D�	 *�'L0T ��lJ�b\U��Г���@��wnk�_��N֊��$ǭ�"�H���+�E��q$�LR�JTo��cO�YR?!��=��:��~�����8��v�	������̈́�����WxU�)��k����$�|�8�m�Iɭo������S,���� k+��IV�d�P�ǐ\���$4K��_�����\j��|����6��'<AǱ�m��p�Ǌ�!dq}!�VTO��W��2ռ#�����]�ޖ`*l��g�����4�H�	=ҷ�cW����LwdŖ+@3i#IDj�������e����W	Mj�(�q�J5F�G�(΍h������G��!�8m�F;[���؊8�I���L�w�R̚��.nO�����&�:y7�|��a$D�s3W�L�#^���kH�0�L���2�{���~uRw��:,<34�Љ��Z���|z�	%i_)�R
�=�f��� �q�,r|���_"�Cb���Cs� '�kV�l�cŵ ���7��G�Y�����R�Ӓ6�%�Wyn=`0(¼��]�Z�z�ވ^�}�����+@��3"%�����Q����w-�Y�U�ܥU;1<o��$�l�B��6���K��	��D�Kz�����qːT�~���䡱S�+�<:H�6؍Q�R��[���8v�Ǣ)c�4��l\�?8R�p|��/��p�O��oq��1d���w,�����c?&��4�B�d�+Ǥ���uUяJ���YG��P���Z3�K̤�JeGl7MG��?���Գ�햇Jto1��1&A9�C��
�$U�wމ':5)t�]2���V&�F{�o����^0a��'����ebl���C�{��	+�M���U���}ݯ������I;����mI��/�0�����\ך����8��9���>ז�����Ӝ�g���,�� ���RઑZ��Y���]��c����E�p��r�aZ�n�����iR��M����p.ktW�w[.Ը����_�&��~g��W�;#e;�\�n�7p�J��Z��	��34����^3R��`(�����主`d�}�:��K��ͷ�V�YYx�n\Qn��}�r/�;�O�F8��D�t�����"~j)���ݑ��~Sy��b_P��f�d"y��"&M�Yޔ����c
y��E�����y�3�3��j����pє}H�ڦ!yM�4H�> ׏����<�%Nݑk��&����֭_u����v����8����6g��:��m�CXA�s��V�*2�RGuIa�G�+1t����n�ǹ����K)yx^~��p�'th��#}��7͕�*=& C�
quq�M��6�[Ϋ�؍F�G�i�`Y�I����x�i�!��7b\��<�Ys�9ޝ�l�ٟX҄Y�bv��;��/�V��c�z-=���p�.��MdC��/���� ����T���.�,��%.��;�S6h��2�y�K����,�I'%˱�O�%�=����ꇌ�_�<3~j=NQ(@J��']�m#P�n�G�>f-�K|�����*�JN���"2�7'�+����$ٳs�q��2r�R>f>[!��~N�4<0}��%b;�r+C����x>��H�����Je�kd��98z�^1pl�jmmB����{	=A��h�|o*�}t&��a�G6���ƫ��Y��V'iݚsn�K7!����F"�s
�X��<ECÅ�;��K��<Tf��zqmn?@��-�vW*O��6����f'M�(�4绸�`�N�`ܡ�O�q�g�|�V&�\���O A��mb@b�;C�%T=���s�	���]�9&�<'��VO�:(�*�f�tL�è�T�	�)�R�@#f�j�lܫ�hQ�SE[MRRcQ�������C�_�-�|��{��������H�W�!
�G�R�F�i=�]�����}�,���G����۱��0�L��q��,��E@ߊ&/j�_UL8a"�2RЮ� s�&(�z$����|�"�E/{'�ş����fæ�� �sm!+a��g=+�_�� �1���Aw�^�1�ćmRL�l@�*��T��4�h�b<�O6'�.���c�����|Ao+`� *�kլ��Tx`���l+mK���*���n��Z
Y�]�X�'�Vy���Lq�f	�Zזr�勿!T�E�ˮܰ��������t�,�D@� W�Dif.;�nsTwb��/�Q����eW5~��u����U�d8A�7=�6Fc�˿�>��b�v����oxg;�ýw��⪥ ���^�596Y�PU��P���|�N�����m�[x^o%�.����QQ�k�ؼ�G,n�qeU�Ǭ�b�K�C�*�mq��a���܏����&�k���c� &��!��v�#��V��p��������ߨ�e+��i�S.���|��\72���fY�?$��H�\�q*��7~�D�6t�ש{��q�����1�Be���q�N�`i`�H0��#�=W����PKyF�Q#  �#  PK  ў,J               101.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG��,ϋ͘��gΜ�]�2�&�gʽ+p�8�֧�����g�xb&�>�&�,riǒ����"m"����Y/���d�P��]N[�uۉ�3Kk�%��<�%X�n$8�1��ڷh���IƢ���"������G��d6��8�xד�,�3WD���X��F��ۃ��Z��V�w^�e��g���F�<�H��n����ﾾ���2�����<���O���iſգy���]J'=�ui,3Xԥ��3/��0�4��XQ����	g/Z���d�����+�=�#%NNX�8�濭�<��
�����j��-�z�g��&�cx��⏏Q��u['�͓-�X�����,�Ek��&��{?g͜���_��ቓ��~p��+�v�e��J����wB�o�CZ�ݳ�%��ہ��y⩏�=b�֬�bu=�/q��W�ە�{�XKn�g�-����&�U�|&�^�W?�&{Q�S���f5�n�E]��K����r�i�?�8,�)Q�)��\��H]ڮx�#��{C��`�lz���}Tv����N]K2%����%�4Dg=�_p�e׳���ז����_%�#�5S�IAC�Qr���2�vDo^��G�S��5����K����.?��A(z�����y����9�$�߅٧,����Jy4���d��wM��H7�bP�w���ס�"�Y�9��lޠ~�)˗�[�@݇�B6��P�u�j�4SN�u�
��fu�v~��k��p>�m���A�����������k�;���ڱ�!4v��6�G-�(x��M PK����  �  PK  ў,J               101.vec��Q�wv�gwwww����݊ݍ�`�؊������v����p·s�;Y��<�) G	JR��)/�d)���(O*R��T�jʏjYDu�5�Em�P�z�O��{�hL�Ҍ洠�]+��z�Ҏ�t�#��Rt��w�;=�I/zӇ�������(d ���2,E��#���b4c�8�3!�Ĭ &铙�T�1��dV*��Y.��s��|��E,fI�b��2}9+X�*V�����Y/7��Mlf[����'v���w��=�e�9�A�C�0G8�1�s����4g8�9�s��\�2W��5�s�����ⶼ�]�q�<������g<�/y��|-߸������G>�/|����K�=R����O�+��w�PK�2oxn  �  PK  ў,J               102.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG��l�6��`S��|~NU��N�	�<Xބ������=�Ar�w~���O��f%�e\tu��XԀ��&:���������I9��+��[�1�aS�'���B�k3r�؋���k��G��,<y'��ݹ>���Μ�g��=�����]����E�㗕vd^�>�S*���K�ffQ�Ƣ��40��|�÷��F^ț<�Q��Or��� Oo���ٔz�����;wO;����v#��b߬v�{j��;|�f�+�� lx���ɷ������g7����r�p�¬.����"80��l���,�"I�Z�{�<�9�qĻ/�zc:�ue��4���:���'Ό�=K�#�GwI�+3� ��/r\��g��2���ܞ�wo9Ӯ|�(�܂^gD���y�'{���ǲ�MT)�z�X��M0��x�T}{g��,�� �oEO�x�R��Po�����.�#�9�����~￶2'm��[��JBƚ�xf��~�޲�
��/�v.�}�u�|�I��K���8gx�a]Ūi��\�Ib����޽Y�x���5���%���V*H�.y]i�Pn��@��+,mz�_��[qp�u���g�=�h��q���װ�6m>����5�
Ӳ�n����~��3G*V�i��Ѽ�~_���^y�����ͷ����gh,�차K�f�?:ѝo��[���t��g�-�V�{���ٝi���S�_n0��_�t����7PKfۭV�  �  PK  ў,J               102.vec�U��P���fpwwwwwwwww����$8�!8��O�e�fe�6mD���+��P�┠dʋRY��z�R��T�"���rQ%���W�:5�I-jS��)?�yn}�iDc�Дf4w�v-�V��miG{:�1��d�Y�BW�ѝ����G����?� 3��)bX����F2�ьa,��
cBV�ILf
S��tf0�n��l}s��|��E,NY,�[�/c9+X�*V����c��z}��f���mlOE��n�����a/������9�O8*�q����9�Y�q�\����U�q����s[��.�����6O�S����s��o��x+��|�������
S|�?���S�����PK�<'�p  �  PK  ў,J               103.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG��l�֭Qݑؖ�����k2�}�$�$�Z��Zb�4��c��c�|���o�ԕ]�&����:����w|�������E�mJ�s�>�����M�Rb%��_֩�ݷe����\'��s��3�>W���~�z����կ������a���GpΓV���v�l{�-�N�b*[v����{���"R��Kii5X%�忌1Y�>����5G��%Iw��<i�����H�D񗥲��IoE}��4��|�#�������,#��������.�O�^��V��m��Z�)�U�d�sa���U�[	�lx�._�ȤԔ�	!�W����/땍w���۫�Z��|9g������	��n��.
�[r%Е���������ʹT@�h�j_K����;Ň������]s�i�����/X��㯫�� ��t�@H�ƋDM]iR�S������ӵ���k>b�u�\$�۵ׇ#�����D��=7���$qŊ��?��1�;���ab�ݺfo6����m������yne����s�O���x�,0J]Ep`�Տe��Y����p<lg�k�v��]S�t������]�WE
��	 PK`�,  g  PK  ў,J               103.vec�e��P��]wwww������݂C��Cp	Οڅ�!��̇I��FdY��rȥy��)�r�d���^�2���@E*�ܨ�ETѫR��Ԡ&��M��u=��^�4��iBS��_s�zKZњ6����Rt��w�]�FwzГ^��������O?�3��bp��C�ag�/4R�b4c�
b\���	Ld���T�1�n��L}���\�1�,LY,�[�/a)�X�
V���α�n����l`#�������f�]��Nv��=�e�mȃ�0G8�1�s����4g8�9�s!ˉ�����U�q�ܴ�%os����>x�#��|�S������?�F�����G>�/��kƷ������)EA���PK7G�s  �  PK  ў,J               104.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG��l�Vͬn�������7���&�}�I֓�ٟ�^�O-t�\��"���E�M4u-d	t����/����w�3f�+���v�=���zUO�{�Ĺ�{R��\W8�����.-�^	�����S��E2�@����%,��v�=>'��ͥp9�����/�J���_�1�ғ)����!뷽��ջ�ZS���������1>���z�{n�=��IF	�/�vT?���w`�Ƣ.�e����sM�q��;�<����3�v��[}����ܒ�w���������%�Ş9\Wi,�q�Kc�7�H���YB���J���������ᱏvG<�;�L#�גY���[Oܕ��o���-.�+mE	E�=��n�ܴz�����~ߙ���4�nw�Ⱥg�]$l+��hO��S��;I��YPѰaQ�̜|��A�U�D�v4�^�z:������ϭfz�8�e�����i�v=���ͺ��Llݭ��z-�_���[��Jh�ޥ5�-�*0o{/���D��'?�����*w}���'��홗|�(�Ţ...�E��iM�͏���3��3%ܠjֵk�3J+��n�|i��e��& PK#k9(!  k  PK  ў,J               104.vec�e�PA�s_���������ݭ�
�؊�؊�`����q�e���}���Ȳ���K��(�(�r�DQR/Ei�P�r��SnT���W�*ըNjR��)/�8��^��4�!�hL���fv�����iC[��>��`�Q�Dg�Еnt�=S�ܯ�އ���?� ;wH�C�ag#�h�06�8���&2��La*Әn7�n�>���a.����"�������`%�X�=�ح�ױ�ld����T���;��.v����c��y�C�G9�qNp�S��g9�y.d9qQ^�2W��5�s��6��m�p�{��y��'<��y�K^�:�o�[��|���)�Fa|+�����)EA���PK`��km  �  PK  ў,J               105.i��eT������ %� ��%8�0tÐJ�tw��Ѝt�t�t
(1�t#�10��֍7�Ž�{^��:����g����5��D�� ڿ<.o,,l�'8��ظ�8xdO	��	�HH���A�tԴ�̼l��L����|�BBB 6q)1I^A!��\����K�O@��)�����z��q�� yh� :11�c? ���'h�-��	6.�?��g ::&Ɠ'������� &����X��f،�d!	�8L2u=�Z�N���>��=����faec���x++�WPT��х��ZXZY�|��s���������92*1)9%5-=#���������������������`phxdtjzf17�����������pzv~qyu}s�����?��"�ǅ������.4t��8c>y��E"��m�J�(�C&��_׃�$�uBn���9��:��������������\� ڿ�a`��&��3��zl�M?+�c���(�m�B��(�>E��b�~o�ᯁ�hK�����ܩ����#�B�����J��=M����y:�q��x��P.�����C���*���Q	�6��W��3NKc�������Q]�	N�9u�M�S��yv���m�"�HƗ7Q�::V�R0w����oA�*fNe�jz�5��5��^�=e��S�'�f���VF@��7�&`�6��V[c�5�&��{K�0N�Y����n"��J/;�՚�#���Hɷ����>�*�<*�*���{��{��9���|�}���Г�[5yc��?��3��VI?�0:^A6�OrN�qD�ǜ��sR^��A�A�Bq���u�a�k��$D�#�|(��˓a){��.cQ�������'��Oc��[+.�#��5uEğup�����@ۍ�Y�W9�p$rO*����|�G�z�u�|��R�{���n�4xz�1�;Th�Q�&]T}�(iK�lM���,��"uJ�C+�l@�u${>tdR���0��V��&M��=�E~��H����șʶk��6���`6�y��SV�Vd8�'^�X�B6K�[�˚�x36|�!�*� cܡ�G�{� +�DA��'�8�u�=�ا=5�F�F[-��ɨ@+�v�uY5��i����g�8��:j#Xzu���� 1r�G@=���D�gW`�2�w���@.���49����y_�R���>�i�FʮC�ٍ-���ɒ�qogaԥ0\��Q!u"�rW�vb��*v��xX�&��+�Z���Dp����#�z/�X�3���bc=-�˺�ɬ�q���ҩ�����<��W%U�m�ɥ|���w�3��k�����������j[�e V|�'�[�@.��Y��1�6�]�V�	���u�����6���\��t���a��+�F}�Lb{�?��ܣ-��&7#.G��1ko�C���IZ�{�W�p�� �i(�BQ2��f����I&����Z��)+���^���Mu������t
���3�=7����RE��pDA�.���G`V7�,�J3�ՠ�ߛ
K�c��jf��A혷( }��=��|��Z� 鋥.Ku<��Z���W��t�X\���/����`�&��7��Y���
�-3��mK���?:"U��7���<\���䒣�Un��m��\n
K�y.�Ϋ���e��Q<�p.mxe�͓ ���a��R�~�cY����a����ʰ��R���/���9�AU��0���Qy��zh�{�\/�����\��u�*^?R�Y� ��G�ӷTjf��&!=)Q���أ��٫�����	�r��;�X�ґ	X6�6pR���-���G|�Ո�2L�IT*�3Q}�ðOe���؆�^�H�����~j�{�?�x��-�O�[*G�7O�R���'��:��mQ��� �Μg11	���N�bz��'��df��F>�I)�!���Ϙ���^���Z���WX��!��kx{��U����.A�C�W�YV���+�P��~z���۷+i���KfϚ�bbZ�F&\z۞L�j�|#a:��}�n����I<����V����{�>���c�T�T,�-6�:jk�g|��bN���8 Ɂ�j����\fFn��`����,�ͫ͘|��&$�������-9�|2;�L�H5%�`ё�zvg��|���O�;��n�+$�o9+6���W�B�=9�w��eǡȏ�MPzVM0����W����7`r����"�!��t,��[�n�oѥ��I��|+ȋ~ԯN�5�K��]A2h_N��������<z x\3,�}@n(w��>�g
]���dĿ�Cs��C�г�C���f��gbMs��;�BYQ�v6Kg���(>YD�:p��0$ge��% ��a<�l*��޲�n>F'�I11�=�O�D�v��+�?1����F2wU�Zx�&r��N�-!�ظ��|·&�w��M�.��p[xZ��u�����ſ<M�\W��7@S�U ���<ˇ���c�ev���gy�ݠ�ʎ$џ��j1�IyS�:��-�z���̆G��sΠ+vL�aoeZ��{V���:�-h��g�ަ����%��l�ZI�Q.�Y�곢B��E "�S0��8(�w�i�MiN5Lw��ơ�0�2���)�,fF��7wC�~���w�Df¡ҋ���&��]�����f9����j�w*�fC�.`{m�ɉ�Y���kyS��$���2���C�=�wCԋ5��{����o�q�)��B�������S~y=�m^��X3u��E���řB��DX�/��L��B-�I,���x�'���3�����]�<X��@������P�~A�K7�"��a�ss1�k8g��=''o���3Y�D��Hm������Y�ѫ�!�R��)E\m��[Ɓ��W��M����k����:���Ĭ~��a,�� z�m�u���}[a�._-�I�=0�h���)	ߊ��G�4�ߩ}�yK�ܬ%v�ƼyYc�>�X{�v��Sܐ�zկO)���&�7����1���aT���@�ک���(�g�����p��A;����60����)���������V���O�{6oޏ��c|���o�+B7j,&2.��BNU��N�%���Fg�4$���؅������⿞���H�᭠�n_��KOB��NŅ��"uY��)�җ����M���]wq���%�nDs�b�Rkw�~3���@�[�S3����A��ɻ�c���7�n��kpjH�|;�����\����X	|#�Uv*kO��b��]�z�&R��g8Z!���(�bp�u�i�y��#P6�q��OBT-Ȗ��ָp~z��O�#�>�q%�Ps�u�I\L���=��ء�B��&�܁��[9UE&5��v��,A�XNɚ�}x~���a *�)5J����R�.�6yZ�~-��?[K'�D��N��,� a���[��,<�lj}�	�N�}�>9B���1ӕJ��j0��^� ��7����?ƶHs�֪�oΠ�	�Ӄ��m�K��&���j��K��Ct�V�4�U\aKRq���:J0f��чͽ[�%p��7�0'ç0�K��P�1�_�w���h���CMBhl%�]�'�J��	R0Hc��ͺ���<8ʕ��p}����9�z�XV�`o^ؕݹ�咋��ޑ6�Ű�nIq�Z^=�[�R�U��Z�q�����
V:��~�a�^����v"2�⍈�6�#���W���6����o�#��x�!�����B/�Л�(g7	[.��v}�E'K��у�X�#�f��xsyw���[h�W����T-\�'��I'C|�c��{[�臨�����x�P��*֒?���ZX�ؑ���\���C �c:/鎆Z�o�0��b�6�1�2�����uP
�giS�w��I��Љf��NA�������N:��f���;B�Ħ�����EWńr\)�MN{���;�-�;U���jۭ[<��γ��V"-	�Km��m���K�Y� �n^,�|����f�˓�u^uVP�*�&5xJK�;jkLQV�H��NNo�]�z�U�'�FÚ�)�u�	��!Fl�Q;G��������W�xk�b������ا���>i��y���\t����<Ę.+�z�z�Qp��:_��_�u@!	�Y���a7�/�y*�]Ԣ�b)���ӉD?��<����.M`��7��E�0Hn��;����2l���gԨ�kwk�ȅ��9�����S����{�9��,ݧ�����
��K�S-+1�7o��(&TrE�д�����GBg��N巾�.W�4��4��a
B��e����1���J�]��ԥ�J҂m�0,-U�7)������x޳�&��IF^#��և'^o���{ĺ�GP`áY�E����(~Zx������&�ʢ�!�qSi2�˳�S%ZR�Â�B�?}��V��J�ل��RMnfF�����zO�Ҝ��ktˤ��@
��E-_�M�YS��3�Z?�t���3���$�g-N('*|y^���.�k9�U�}]�F�uIZ�涣��o����R#l��u߲8��[p�&̪�����7�=5j�{I�*8D43L[݁yE��jV�F]{\$r�)%�(q�bAt>�?�qX��˭�Y����4z�6Ԃx���\�_+�l*�Ƅt���̺��-><���;|y
%p'��0�e9k!k�^�f\o�̒���R���m�W��S�9w7z�)S�/Zm�P�y��!�=�����ͻ���s�*�_��YtK��b�9��>n��ok-0��-���_�;%B��	ƃ��>�Q-���3�
�4�\6u�:���.�"i��l�6eNa�~��v��{b9�|�u.��������~oj�?������m��&i*4�p����u+vĕ�W����_�\I1���02%�n�ck2�={���P��f���}�����y=A.&
-�����R�> Mi���n"#GI�&�`��
�v^�����P���:~����F�F��JU��7����.�S�E!�g��!�O[��P�����/W<��s����ЦP��c3ڇ}㭋�����9M�	��߯J��m�R�˭A])����,gN����}�3�f�>mR��i�_�Nݧ��?.�QX�=�y��sӣ"1.p\17��OU_���I��<늙�ͼ�0�M$/0�->g�h��P@m�"�V� ]�Y��K��΀A�W���ʝW�
7�"�Rd�)٬�E�����q#0���y�!��t�cB���H��v��<�bS���3���S�����猈u�*����Z�դ�@�j��2>���t��~��G�!pg�-��!9�L�P[~�j�uHd3����=^ߏh���7\���q�z��
˃���ͯ��H�Dyʇ��]F�V�q� ħz�6�D����գ���l��7[�^�~�U�!��#���t'�$X��ͿY_r�.��M5-l�t�Y�0z�*���۰���fV�$K<+~k�Nռ��n�ɶ=�,��"V������F�;�$(u���J�,����m$5q�̰��n=�[2<�J0I�ŝ����G@�D���eP�-��\n��@WIT�ݛUWs�,Gl%՛���8�/8�ήr2���sq#�M.�7+&��U��=ܞvm4�������#�j��>�w�3���',�A&����;;%!rI���f��D~$�}����l6����'��CV��q��gЂ0�@�����`e�6�.�N���B�I�C䒪�<Cw�$��/��1��l�Hp�0��E�9�f�nS��Q���B�iN�R�l��"F�g������@���~F@"��-rA�3�Y\'F@�����R�'����#&_�]x ��Ր��3/˚Q�թAm:���o�y
�����]��.��w�[,��1��r��B�uS~��ž������M���q[���z\�@��G��<�Bȿ�']0�>�@��gg-Hh��y��Dc����^!�z�~_9[ƾ���.�$�h�ԒP����%�fT����^n���N��E{�(F(����j�������v	Y�t�X��Ѧ�C�7�֣"?̹֮���c�Z��*0Q�/q�:�IS�/���[��H��KDYߺƺ�_�x�/������!��2�i�`|��s�<�����|�K������>J�Q��	6�S�{�K�EO�FP�<��:Ͱ��3f9GT*K��*�k�����VOd�����1����3n�{L���L�D��A�/�&|v3��[]����[�!��Ee���ae�H��C[�e�~������p�rL���N�p�G�`��x�/�t����lՎ6.p���ڍ�@6��X`T�!����/��CMp��
�*܉�̞�Y�����?����_�"�*�z��Ѽ(�����oi�_��w!�(H�p!tj�f�zH�\$�������R|���m��o�[��.��߾7xmM>�`UO��p��2�[��?}��E�����s׏C�(���8��B�N=�rc�Jbs5b��y�m����_��qS���y��c�F��t�}��~�	�R���*	��`�fJ���D<9����^x���d����]~���sd!���	�}�L��^�d�{�|���B��~��t�p6�o�?���9~��J�8�r#*+�DmP��8�� u�-����U������~);b� ʻ�0|�"73���:Z��Ɩ;UY��� ę��2|�������gZ�n�(���r��5N&�1v)w�R�5�ث�y�?��������O���n��;geUfN�	B��D)���W�yӫ����Z�֩$y릑��2�K�1J�����Y��cU&�ku�PIK�q	��`%O܍%y]R!/Y����V���!��0��������z��6s:���I�o��B�r�)K&&̭:�D�ޮ�͜k�8��@a
�Չ�f�|͋�����l�|{�����G�z G�eC��e��W0�ow���Q{��~���&��{��w�ō�@�L��W��}EIc��o��m骫f��NrKv�e�ɤ�CXPS~ꎅ� ��*��7���N���m׸����p*c�Y����������H��t3_�g�s�լm�!n��ު]��U�y���P��	�&=��E����T�3�����/ΰ�J�{&M�F��k��'.�
����D��/Z����2۝�k%4�A���o}�����7�c Me�o�V�|�
�ݿ(w$�񺱸��Ϲo�|t=�}}���w�Id,����M�J�/�B������{��T��z����D;���t�m�~e����Fj^Re<����~�j%�o[�q��h�G�z�ƭ�i�YVZu}n�:�P=��D��ُmyb��X~��_���6h��\�m8�V�	�ï�K��s{d�n<{���OWB��@,�]E4K"*�Z��0nD8��9�%(�#�s�fd�(&H���9�Z�#�$"I*B�EC��+���
ɾ�#@��܌CT�\�cA�=���¼btï��-2�|���n��r`�10�]���P_��\ԩ/0��G�+7e[��8���I`�Ti��2�"�گ+	��~�Ϋ����;��Lv3�O	�^f�Gza���7�ϰ�@�ew`Mw4Zħ�I5�0��~�� �K�$�E�ST�Ϸ���P��r�MWQ=��,�ݙ���A�C~S�׿^�qO�/��G��O���r�z�B5i�u��>��p�+U{;u4W�^�Aq��U0�Z��h�@�����z��"L������HG���k�A���Џ8�a�Eo$���&O�%��d��eLW��Z�b7UQ5@2�7o�w��HK�=������%���2Ę�N"dY�!�k�璾��S^"k #�˄��@	=q���9�	Fq�E�Wf;ez�g
�Ϝ��nD��~�;��ﹴE<��ѩ��R�k+\Vzzj�!�[�����;|XSz�bu�p.0�2�;�S{MHExt|Ů*�,��W���t5`ju��'@�`�[@����G��Q�Cˑ|ܮ����~�v��Zy�zZ���.���8�ݼVw3��W
�◣:�
��6�ȺŎ������J�0(Q��>Q�qn��kp�a���D���Л]��i�*���a3�M��anFa*څ�`�fibX�2x�"'�������,�1�_`�0�z˓��cQ�/�,GW����Tާ����%$Azy*�ETz�'g�<���P���^ÅT���������<��N��I�(-r���|H�~x4���n�J������ *�\tPu�2�������W'�Ӵ�V��|Y),P���豮����Ni�{*%�H|c[�b�	�RBw�������wf�%��UE��\�#��{�k9S
aH��:���1<Q$f�0�~��$�Բm��8 ���?�܅gi��n�l�KّP���R�M��j�V,S�w����Zn�*��;�x��ϴO�$����g�L�B��(߄������LJ�5���T������b0b{��44��v�O�E�|��ҟS�M�ߐ�ġpf�\���0f� ��L�h*����+�Fei٨"�Nor:)�gXN#��Ei��ҁ�)�u�W��=t�8�w^��'�v��=�K�[n� �����'��gU�)\��	fs[֋�u��*�"�6�Rx>����O-���ysD	�t�2��5 ���S��m�M̸
')�qi?.�PK��*�"  �#  PK  ў,J               106.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG���o�f��A��'i~0�K����®���k��~}��E^My��g��0�
��{Vy��.��@Wz✬�{��3sm�S����;�c٫�����t6��w����~Ϧ�+;ui,SXԥ��3/����wdW7�����K{�����6V�m���W�|vr^(���u�Z`{Nե��/�)�έh_'���Ɠ�*�3\J	�7����ܯJ�'<��ۺ�����=O7�_�"��eJ�k �H�.,k����ʙR=ǜD�N��gS��c�J�ױ�6׳��9��U��v�I�z��2�&��,�º��IB���A�����N��W��կ\w��TIج9�"��e���=�ب\})��zZƢ�d.�E���Gӛ��v��k-��r�q]V�����M�W,��\�,;Stѧ<Ղ1����.�'"�kVfF��+�]E�LnV�C�s�T�ĀV�e�"O�����=t�$�Ptª�<uS�n�g�t#���^����@W<�q룟{������`�J��l��l[t:|kѩ�y{V�_���A����o�K��6����'`W^\����j��g�/(�U<�gNx�����*ޗ�Zn�#�ZS��_��'6�2ޥw��q�9�B�'�\	te���{|+e��,�q���`]��-�/�j���/�t|��c]":-�a��Nb��� PKl%Qb  �  PK  ў,J               106.vec��a�w�k��ε��[��vWl[l�Vl�V��Swe|dx8�����LD���+C�d)Ei�P6�D�$��^��T�2U�J5��yQî�^��ԡ.��O
�l4��Fzc�Дf4�-i�F��k�����@G:љ.��j�M�Nzҋ���/��W����� 3��c�݈$#�Q�fc�x&01�Ť$?&�S��4�3���b������1�,d�Y�R�er9+X�*V����K�Xo�A��&6���lc;;Ғ�i�K�����"�������9�Q�q����9�Y�q�\L2qI^�
W��unp�[6���r��<�!�x�>�Oy�s^�W����M�7��w����g�/�k��-r�=W?��I.~������PK쨊�r  �  PK  ў,J               107.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG�c�kw����T�Wjb�X�d�b�,�e���JZ����si̓{�l�<h�ظ�Hzμ��.m���E]����o^e8s��� ���M�Ź);��=���?ړm���ӣ���;��+�v�3/n�W���dF�J����=�b���I�mc�*2n�y}�C�fY������zlXԥ��3/���R�^ذx�C�w���i��]���Zs��.m4z�/�8{��3�~��b���Rg��»6=���x��������Ѯ��s_ʹ�%R�㺩��<������L	t�`	t��e�6LO���~6Y�l����{&�9w���z��]���O?�|�i�gsL��S�����uOM5l�c*�d����j�.���po�ڎ��3��\w�ȵ��}Vt�2r���}�_�>�,�{˻b9��=��X4ӑ@�b�ޡ�����ɕ;B���<�����O���e��h�8��Tgc�É�����c�^�ݥ�������좫�X�@(Q��(�o�V�;�	��'��˯-�������s�?�oP�r���{���9Nwg��z*yضw�=��u�P+���'�L���{�v=��;�����	�sr�f��xWnU��?C�]%�U��ӗ9��?�3�w«��	���hJ8y����On_��~��$���x��ϧ�,���&�Y�nɬ���)W]Y�Œ����ٝ�D�nު.`��:l���YNyo�ݛ��z�K�B��� PK��1�  �  PK  ў,J               107.vec��Q�o��������������[��Vl�Vl�?u���6sf"�,�_���%)Eiʤ�(�E���S��T�2U�J�T��j�5�Em�P�zԧA�EC�6�ӄ�4�9-hI����]�-�hO:҉�t�v�����'��M��/E��~�1��a(�n7"��H}��X�1�	LL��d7Y��T�1��d�������1�,d�Y�R�er9+X�*V����KY��۠od���V����8v���w����c?8�!s���8'8�)Ns����<�ȥ� .�+\�׹�M�-y�掼�=��<�1O|����y�K^�7�͊�|�>��|�+�"���Ǐ|>~꿲|�����PK�X�k  �  PK  ў,J               108.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG�c��.�����?��5k�y�bɄ�����G]�z:w	����uF\g�]��d~�mj۳kӌ2u%qi,j�'6+�I�I��R�%׵cK_�(�f3�ͩ��O���ĥ��7+��D�
/T{�R���c���v\�H��}Q�:=|��Bw��S�?���?��;��+��4v�" �U�f��Ux0{��2תM���Ә���~m�ܸk��}&?��|����#է7~_�ȫb�j0sQ�_b��wE�?;�ɕ�}�̪��ۺ�w�$��_6=w��Q�uɚ�˦wj9����U$��5ۜ�|��%��Og��u�ɯ-�$s"{�5�W#�.�,�W��f�����|�0+��竘E]�=���ᗦ�_,�2��S��@ቓ��c�zN=�s��Ѥ��.��uu��m�������lt	� d����[v��'�
n������e��Y��^�Qm���-$����Ƭ=2��{J ��e�:�恜,�/ @Xz���$���'�훮+ݯ�������3ĂN0}}?�m���_�lS�;*q6,��`���ݏ�gW���y�*�W�=_�[fS�K��U�w��m�c�o͞i�k�Q���-�#����;5�����[7�D֚�:����TU�w��s��+n��I�
��n�+�3�f�ӏ������M�V!����������U~�n���v��c�՝����l��]�҆W��o PK�X�$�  �  PK  ў,J               108.vec���7��g��kww���]��]`�؊�؊�`����{.���H����(��<�(M�f�(�D��+P�JQ�*T�ZV�ݫ�פ��C]�Q�Y>�5ҋiL�Ҍ洠e�E+��z�Ҏ�t�#���^��z7�Ӄ���7}�E�K��_@	�`�0�avÓ���d��X�1�	Yݛ�Of
S��tf0�YY����s��|��E,f��R���`%�X�ֺ��n����lb3[��6���v;�]�f{��~p�C�G9�qNp�S��g9�y.p1��%y�+\�׹�Mn�7���r��<�!�xl�D>��y�K^�7��x+��|�������[��=M��3I���ݟ��PKEB�%j  �  PK  ў,J               109.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK]EG�c�,MO���zB��hIF���S�$����ߝ]=�K[���Z��2��.D9�n��X"o��)���Ϡ����4]E�7�9w�8$�y%����k;�^��Hq?â�����U;���RN�}�혽:�m�2�����ϙv�d�lxsl/�Q�MY�^+B<&��)�Yai�����W~^r>�٬��E]��p�[#H�i�1bT�k�����%�~]/_;crDA�i@�K�٣��W�_��\���r�J�}�6�',��z�Lz�ͪ'�_־^=� SU�a�fc��
�
ⒿB~Q]ԥuD$Е.�:;� �.HMD\���O�GN+�����1_�j��^Jw��O���rƖs�l�>��"�>�r�������g�2?yj�9�g;U��L�{��NewS�Wdbij�1[�ߤ��}z���K��QS��&<�o�Q���8�U�\�ڙ��Ǭ=y����y��#��z*��nJNu���Ƶ��w�4�3�Gef�\{zKc���R���g�7Ϙ!zS�/kQ���k��Eo�]��q��`�W��ݯ��5���Ů"!��-�=29K�l����D�5B�*���M?�"/x�������U��NR��"*u��{�T^+�.��׾.�j�ܠ����y�����r�|��y������z�����	�;����yOw�[����F��,�EM��!g�y���K�<��~���.:1�N9�^�I���3.�ʶ�^GV)���	 PK�СF�  �  PK  ў,J               109.vec��Q�o�{��������V��.�[l�Vl�V��S=.{3l���,��O����)A�T����z�R��T�"��������ըNjR��ԡn�E=��z҈�4�)�h�R��k���5mhK;�Ӂ���d�Y�BW�ѝ���SD�,}�~�g �`�0�nXV���d��X�1>�c��&ꓘ��2���`f�b��l}s��|��E,�Y"����`%�X͚�7�ڭ�׳��lb3[��6߶�n���]�f{��~p�C�G9�qNp�S��g9�y.�㢼�e�p�k\�7��[�6w��=��<�y,��g<�/y���O��oy�����G>�/��k��[>��Y>~�_����PKC�UXk  �  PK  ў,J               110.i��uTN���� ��,�����"���� ��,ݰ��(-%�J#Hw/H�tI����{�����{��c�=s�3w�����[�+�+�p  8�p7�<��'��{H@@@H����1	�G�4�Td�h�����L��L,�z�g"Ϲ��_�|	���
H�
��oBBB�G� � 3=���g�kP<đ� qX (p�8w] ��9�p�����< ���<$$zt�"<����pq���~ .%3�>����A��!��;�5ƏYM]�	��<�в�s<{��RHX**&�ZN^���������o`���������������'$4,<"2*:)�SJjZzFf^~Aᷢ�Қ�:ԏ��Ʀ_�]�=�}��S����s�k�6��wv�����_\^]��ǅ ��o�䢸�z���%�����x����2���X�>~��[�A�8�6u'z��r���h����X��/����� �@���) 0�߽�0��ٙ�F"�Z����$Y���d�v���(�g�+���°�:[g��5묷x$�����H��U�]���O����S�M��H���Bc�2�tَ�G�xn5����>H��Ņw� v��R�=��z5u�%9?�n6Fү_�����rQRXt;%�3L�{�[U�bP/�����0(���k���
\y���_@���]$��E�ޱ�����jz�A�O�S���#���.DW�;�:�]��z�������'	�<*���ץ2�hƠyj�^�DR@��ݩu�\��$��!V�h���;@����X�n����.��%�Ąa)�7O1L��rr�-�+K�4[=���:���Qx��kOJ�M�ݬ�B��Nzv\�s����{��Q骅�|�#1a)d��y����w%�?�4�&�e`ݣ�*��v�̪_7 ��R��v7��� 8��
��-���VEĝC	�{�5�Ϙ���s�g8Rr�f�nBo'��@��S�%�{���s1�Ո����2G�r�S%E�oʸ�0{�
6�>A�E�����R�5.E�f�[�y�x,�Ӭ�~*;�%� �l�l������ԏ|�0��4&�; ��0S��["(�'σG^�m�
�
�B�DH����a�7OL=ԇ\�?���\��Hs����i}�7�y������U��M�35Ξ��`�?�V-7Gl�Z�G���P���F�~¹��{��FC��rK^_�X�jԎ�U�tֵ�H���c��2[�Z�:Ω]�!
d��R%�8�>mj�0��{���gZ��;o�����V\n>W�47�<%�Y>����&��Z��6��a��Mz�r�M_�C��j�o�2��mM������i�P�}[۰Q%^��Q%e��������e�!�����(�*Q���(�Ϟ�r&��fL��]��ZLD���i8�1F�����h��&\r�Y�獺�+'���n����ZGNL0)��1����R�ۈ^�s���rz�r.G�y�;����V_��Xԣ�|ǧHc�hL��w�J0�Zt,�)��.4�D���y�R)�y���$�zX�8���"n��O�3�:�3�r��tMN������ W_Ο}K�[cd���v/\��Gϛ���>����|ݺ]]�m3D�F+��WY`�
uOu�h	�ي)�IhW������\%�GҮ���G�Y�bcMj�b��٦��G��yn~��H�� '2?�;��������%��߫�lzޖ+��!@*rcQ��9��ۣ]<�R9�g�	]���OC8��ߨG=���a���uz>JyY�&������vڜ�qD�򃴶����Y)KvN����e�5l] �M�b�}W�Ɓ���y{~u���>�@�[�x
���-w��.o��~���^e檐�>_Z��v�VW�4��8޻ґ��
��7`d��?=�#u ��p+W��وX*�zM�c��wE�➻���H��+��-Tj����"i���v�>�@�J����v�~a�f�/�[.��1,%��N�t��j�9�����哹{FX��@="����˨z��k���� O�+k�
qycӃ,��y�Q=����S
5bX��T�3��rafI~А�)�0"G��n�(��*��Q/������F��k�����^�"�iX��J�-�Ĳ�s9���9����g�͏���A�G���8��ky3E'�y��Ѱ��V������H�Dg�v/���V��m{�F�Gf+P=��I���k�0����U�\&��W<��S�d��S��es�5
.I��,�W�S���>��|iI�#��N�6kqwhAp~����_��4]6;�_%j��c�,=1U�G�	���L�%w\�	���׋��&l�޴'q�S��ʢ�0����"ݪ��h�!��o쯜�vR�����i�DY��iG�	c�ʏ�{sF��>����&�v�jB�ŀ�^��'�O鄤���|��@B��t�IlN#_Ǟ�K��t�G�M�qL	j��D���l ��yidJ�m?�����}tu���8E��iȀ�����F`�:x���+�6�T�x�p��,6��U��YQ>��Zl�+t&�Д�8�(z��#%´6Kݾ�̈��K������W�<篂Fь8YC966�"`Q��6�@Ea��G�_��녚�jm�DA��{�Y�/�F������?��Zǋh��uo'��~W��$t�ܺt���@�L�f���/
P����������5T[���8���G�o�O�c:R����>ڴ���
�]Oy��PC�Y\���͚y��ꎳ"� E�y_-�$E�ioʘL����A@������a,����ה���1,��ןL�e�����n�U�
�ƕ�ƚ]�-��j&��AP'G�NM�WN�Њ]�t`�V��Et�������Z�yN��_>�Za�R�i�����Y�-�N�eR]�����
��y�!����_�b�H��:�\z���.��/�Z�s��٠� v�LU�"|u9�����*�	��6,Hz�5(Ы£1�=�T~D��$�9�-�W��;%��U�.�\��;�$�	�_ \;]��2X�4��L����|'%z�w+��T��RQ]p���|e4���Z�A�@�ߋ�`Ư�v��� ���;G��2��{�<T�=�m��"����=m{�-�=��P����@�=L)6=�����!��\��k��޳
��A���b����)$I� /H��|e����A�wLU��$,u���(�8��U��0OY���@���+,���)g��Njv�&	�5��D��
]�d����iKͲE�rU�}�^"��Z�c�ܬ�Q�k��KK����i��=J�����3v��L�U�����{Yf�X�}���_�8�n^�PiJ��+�I&�K1�a6����~�sM�0�*���[��±:\k��/2=� ^S��Gϰ&01��f�_��+�JE��$:�	�娫��A���O��k{ϿA	�����Ѱfn���Z���� �~;���1��]]���vͧR�fX��ER�}&�L�K��L���wN��d&/v�t%��фD�c.�C�2�P�e� �'�	���ݥt1�϶z�c�+U'�BQ��9�*fc�5�P�@S6�"���=���=�w�������l&	�q~�#���K`)_�O��޳��fr���֯ف�Ǩ�gqq��H�p�چ;-בL�̣�����|]8QXW�J����`�������X�1���e��|��
�-��f�T���_%>l�m	��ygX�����'4`X?�lв����2_kv���Wc�Y���*N%;/M�(�������W|���1���Ђ8�>��a'�c��
�>Jp!<[��V��x����F�$O������MU&9QK�z��z]��2{?D�=M<��9��KJ	�u�ZV�{KD��J���F����]@q*��
��!�rq���@���n E�Ԑa�Ʉ��H`}�w��gZ�|Np�\�Ш��\*��:�#�GxCtn��x�ͣvT�M�fq��-��؎�7c�O *N�.a�'��"�sh��$��b ���	��l��7��9��F�V�v�G��z��ȓ��N��ur�/{]��'����N��_ʭ�MP�S;Kt��eSEF<�Z��)2�{�b���d�}A�߻2m�����EM����?~���I
GD~�E.��al��b��d�%��G��x�̴�AYӈ��B&J��u!��J*�ٙ��)vtm�a�"o� ���k�&�!^�ΏdW�\��4�#� �������!�!�:�r�h��|�16#?�&�n�-V�z��P��*��&���hYl����9E�d� ޅ�3��9�r�w�:�s�P�#5S-�]�gŻ�d��޻���������~l��9�7�ݚӶ�N�w\P=9_�`#߭R����i���9 �	�s�+֓���B'��� �T�U�RM�]B���^�X
Z��ʱn[\�Tj���������9��;�3p;���R�f�5�^Y?�]�7�UF�XL���نBII�t1�����Tÿ�g��ŕO�qo4�̻�%���o��;~V����o<T��L���@�A���rb�Q�{*�j��� ��qi����>#�7ʋ����� +��&֊�������!�\
�Y���߼z�	�?���d7�P�Ó��ힺ����G��q�Yo>�q�������T5�+C�(��g_[��<��rߵ�.*����(���,g���l8�4$�z�1�#ZAv��� �6~8�C~Yw�*T�i�C8)�p/���1�Ҿ����J��Xz����UK����7 �.o�����̸k�n��)^Y��ɭ��Br6R�T9��T����x�i'��^�d�|)A����I�L����*�c�S�{�����$᎝�������2C�w�}O���� �r�븨��Z�������l�k���U� �!R��|�Iln�<w��G(|�rä�^��&��ܛFJ�̑��0iYTh�U�E�1#��&)j�b٫^^Z���N"
e��O��Hc�J����R@s*=�� ���+����	���-��!�
������}�/�e�n!� ry��n[�~�����~�<�3��H��GC�M��%���2�����NE��v.�N��	DN�-�{�����tv���^�u�)���˛)Rd��Ӕ�A�=uɥԚb��{��</'4�:�]3�q֎�B!�_�:����tok�9b�dF�ڊJ����>M��T���A���bq��@d��o��O�?˟�W����U�g�"����l6|�< �BS'���Ǹ*:�j�%���W�Uh{̋P���i��Es�%�I�Wc�5�P8���x�!AHv�؍�M:��9�ԝ��@�(M�F���xɒ_Q�T-�����δA��<J�H�e2x�O���ٔ�=1�Hf��!5%���[�K<> ��+��f��\MS�����2ɟ�E��r|�7�����w�=+h�����N���ߖ��}��a�w0S~�7l}ӻ������cYߊݒ
�����!�D���=K��	�\
*l]9��'%%U;��J�-���m��.>��rO�!&u#_v<\f�f��:=a�c]�xhއE��y;�&J��'���
o�
��%	V�+)ݽ$~d����6t��f;*Ҵތ��&P���Wh�4W���=�Ww ��kZ1C�&d����>{W�D�)�,YQ��N9����#w�c5��	~u_G��6ǭ��r���-�L���4z�'O8��w�.�jr�O�V3�L@ 5[�b��uOl�r%yb)�g��$���c뚨�Ģ�}�۰�����1�5�/�~��艶�2��|��%^�MT��ʁ�\{��aQ�DQ}���k�������9��ZQ	��p̩
�m�xΰ�/V�FR0�"����=��u5��]&l�1C��Ց�����eJ1���;!8���TD�*�{�T4�a�B>����x��P)�/�}�eWN��Eq�/���:_����m���?�R�}�7�!-�22Ǎ���,ۖ������kBDV[�؂?nT!Z��J��U�+-�]�;��.��ڙ��L�
��] �hF��m�����ky��p	�<����#ar�Į ���x<o�ߔL�x��f�lg��T��76H��Ee�5�����7���z&{��j�S�Va��<���i��ǝŃk�%*�� ��W�5Z��i�7,rnP�6$lF��y�1�f�pr��Y�ވ���f�hKh��l\�X޴1��Lm,Ʀ�3�o���0$ٸpz�3wԦ�ԁ"h�K/80�d�Z�wpp	wn��Y��\\�6���ܨ�<�Ʀ��D�z�Ò6O��tӘ_p�d���� �j[��G�K�@�����Q��+pz�k��/9�� ��j�r�z��M����dyR0y\�mPw`"U�m���6?u���d�(�����4����L�. }Du��1�%^C�͓c�#$�A3�T����G;q�����JH^Sf��/O� ��G%}�ͥ�	�-�~�k{�y�V��'�8-&	�w I��Sy���=��2��?	u|.C
��]��寕���n1��@^�ć�'�#0*4��ȉ���w ڮ��]���\�M��T(������:�~�����&�C8��B�OhL*� ��f�u���)5:��M}W`9��䗍�~���M�(���z��u|��t"��ϴN�[~k=���T����ږj��*��̆��}�[:�����-*��T��*�`,;
��b3���~6��I�b31ad�2[�Gg>%��y�N?�N�7���4hN:kx'�����Մ1����m_}Q�ھ�sc�m����9|"�:q���μ;�V����i���?�,��떁Ż*�J��䵸y��@�P �nO=T(��QnQ��F�<�sq$����X-1��Ԏh�1�f�DpV��DL:a-ʴ##����r����.!��z+3�Ų�d)�a��O6q���;�3@W���R�O4��Z��E|�v뺈�\��W�jgt��:<�GE=��G��7�������;�����������'v�E&�إ�9S�%	��ۜ��"��ª��&SJv�E�����XJ+"���;�C����U���<����G���'
?Y��������)E�b��gC*���w_Q$$� �u�N)�EW�W<"�����/_#�����w �� wzʒ�?G;���1��t7��~�u0'�I�V��)d�'r+K� ��d�'|$�R-@�9ҸC�nW\�Y�VHҩGG�uh���]�L�����0A��.�͈���U����e,X�T�=4���Lp^��0�2v�tV.�7�ʃ,u������p��[�ͼpX�+5;�Z^��(/im���e�~V�7�o��4�?6Ŝ�w^S�^���=�m���MSZͬf�P��¼�q0%7n;�?�~Z��:ʪ!���d������U)�e�`���	��w/�>}<�gR�5�K������s'��2��N
�=��FJj=�Cp6'����Pg�,1�֐�`����3+z5$���s��Z�d[��p�^5Z�Y��r@�3G�f�����t�oi�t�NWpW��H��|W}*]�^�P���o�� W|��i�����JR�?��
��'9���K�1�k��D.W��[�u	m��������s%��쪅*�Bɼ�&K���|m����b�N��R +x��Lĝ�<L,�*ٌ<��8a�!?hz'�/��8��_��獸̛�]�����4_h����	잁'j�y��8������d"^>xv��A��Op��Ó�3[����k�D���Yw��s��&���?e���+�AR$f{�oWwT����{!*A��p���dV�l�9cX!�cA���օcQ�^ܴL� ���46�FEVdB3Z�O��������eO4�UG�4��j��~�vZB.Þ�OJn��1e���fY�,(�����6����|z�=/��rAw '�?�-�U��/�b�9}�>�&�;?ɶ�6����٥�p��3c��\|Н^�Ǘ�*��fw *M�n�F�,���H��Zm���Z�势��r��S�Xx�tJ�M?����V��ͧ��1�5���`�7Z�=�*�f�K��9.�e7�ui��_���H���o����?����H�?�@�ۿ���O=�^�v������y(��tV��W?W�����u�m�}�g�x)��($أ
y_���
5�o�֒�݅�k�\tf�[,�׋֍�W�~VT���%�ܝ7�>TK�*t�Le�Wt�~�h �:!���-M�N_j^F���&�7R��m4ɵ�M3���%n]�ձ�/ڟ���O���艪d���ܾ�9-�4���]�u������ʵ7/f8��>� J���f��U�^����@Y[��>R1죏�I_Ԉ��/қ��̴z�trh&��h54
�0�9��u�j�Bho�2 On�a3��9��Aκ�Kb��]�u����3K���w?c�,����&�/ƣJMY�ͺ�/U��?V��Ã�"��&wT���W��J4��D!w sjPT�����"'tN�@g4���z�F�ɃU�T�޾������#��ʖǩ9�M2<��%�iz�����'�׺Vw�'dJ-�N�^���`�g���O�%0#��O���8��kv���u<m��ٕ�}��q�U���[	�P��UT3�9
%Ҟ�/�]־Fx���?I�6������PK#��#  �#  PK  ў,J               111.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK��4����f�7>}�^x@6;��,~��E�s��z{We9;���������}��Dϥ��:��N�?�Q���ճ��]E��V�j{^�ݴ@�'\�/{��)w$�0r;���٦n����5�~�Vd��ǽ�݄w�������,��������ݟk��X��Ϻ��W8�M�<W�?�ݪJgEX�`Y�uy~�K#f�ܯW����ޯ�G��,u�~b��$G������X�����lV���'ω�O��p�˺����mU)����S}����'��T^����0�Kc��Ƣ.\�U��ݙ[�,�b�����Ƅ4�\~�����:�ă�!��.���IK�5K�|�NW� F��}�M�eKU�*��*�'�X��fs��m�*�#��{�X�#�Ιl���\٥��vrŢ�d.�E���z1�7�'�������cwn
1��4�����Qm�n�V�-����Kr�y2�S��;�]E�t��_�����if}N�j�3p=��^~m�<�)��620�Z�gh�zr(tc�n+i��ʾ�?�����Oc����u��n�w;B�ݶ"��h㪦]S^E��{#���.d�DYd�g�j#�T��=�v�&�?h��Oi�h����w���zv�r/���2��k���w����Q*_|�,X��+#q������0�]q.I����*�9��2�^֘��W�NYia�'mϮ����q쑟f���;ہ���ef�����9*qh�T�K_�G��u���}9k�2�w�Z�*��& PK����    PK  ў,J               111.vec�e�VQ��:3vwww����]��]`�؊��
�`���q�K���lΗs#�,���O%)Eiʤ�(kWN/O*R��T�*�R~T���פ��C]�Q�� �5�ӄ�4�9-hI����]�-�hO:҉�tq_�,��ޝ����C_����Y~�R� 3��cx*�Yq��G1�1�e��Ĕ�IYAL֧0�iLg3�������<泀�,b1KXj�L.g+Y�jְ�u�o��۠od���V����(v���w����c?8�!s���8'8�)Ns����<�ȥ,/.�+\�׹�Mnq�ޑw��}�G<��S����%�x����|�#�����"�FQ|�\|���G�������۟H� PK��;um  �  PK  ў,J               112.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK��4��ǜd��-�|���M�nG��~}"���{���M�;ؿ���=�*}V���j-�����X��E%lbZ1崅D����%d�/M�̹���D7ǰ�^�޹�(Y�kß��Oc�=�	9�R�Ţ�EN<�{��>�˴�'N������n_��Ӿ.��}��/�˟������R��y���#�2Jܑ�y��8�����3�3}�3R���6���,���fwY���y{/��]E�ui���˯%N-�d��zr�*[���v町�_Ǯ�p�w崉ʑ'��N��g�z��\��u��O�ַJ����{���3���)�a�6������L'ZO�sϪI"�p�m��"�a��"80�������d���LM<q��qLr�9r�v�V�X��uj�i���j;
����r'�������}�m��d�݁E!̷��_v=a80q����t/���n[�����~nqПm��;��6�u	0 l��ӭW�����q'�	�
j��j��U�H�M/�tH`�C�	�u�'u�}s��f��*"��f�ȋ��*�m�J-��׳���ז���?���w�τ⋬Ek��_[��uw����f��<ۣ%���M��������(�I�F��?�՞y�L�-�J����_槕�.d�+B���?kZԙ.~G�>u����:���G�W�]{�' ��g@�c�z����_Ԭ��^r����>�E&uY�N����n��[-��[���s��j{����.�G�+c�/�"P8��z����z=_-�U��z0�p�s�NE�ӏ���9-	ek�._}>�qĮi�L�S67�x�l�V���� PKV����  "  PK  ў,J               112.vec��Q�o��������������V�[l�Vl[��SW9.{3l���DdY��J���<%)Eiʤ\��+����De�P�j�(����kR��ԡ.��O����v���4�)�hNZ�*�hm�FoK;�Ӂ�t�3]<�k�M�Nzҋ���/�RD�,�3��a(���ƈ,#�Q�fc�x&01b��d}
S��tf0�Y�NY̱���c>X�"���6��rV��U�fkY����m�7���la+�����r���^�����9�Q�q����9�Y�q�\t���e�p�k\�7���ݖw��=����G�o�D>��y�K^ټ�ox�;g�^~�#��̗�_��
��)~�_����PK)z�h  �  PK  ў,J               113.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK��4���yuS�M�}�^�� ��Ϭ��4B�&O�z{��«��*+D��g��V��J
���X�b¢.<���i�ٶr�}�6���W�P۝�u����.�Q�RE���u��~�f:,�����\��j�Ԅ�}n�V���NH�7���[�:��̻6��
��V��Jl��1�b^QJU�f��:�²n��&�:�t����tKu�;�O���~�?���y��J��=��%��������j6ǘ��I�)�>�zj�9�og�'=yU!�+���=������N��ce��l��"�a��"80������Y�&\��~�Z>W�?s]�ќ�9�S����^�e�N��=O�\g�Z�.#��N�.?���ޕ�i��au��c����1��W>��w�mߡp木ྺ=�3D=[�3wB����"Uk3_W�� <N;���}�^E�l��jw$\�T�Q����ϱ���{Ĵ�N�{����죲�ďd �u�F>lZ�k��:z����OƜ�}�u��#�=KW���δ��K���7ǹ��Y{��B��2�Y'���u��YU�[��t���wϭXzE�_Y���f��D~�yk����̌W�[���<�6ӗ�;��������\��o���N���;S�OO��Zk�,�4In�wR��WR�s6Wx}}<]bbQ�#����?�ύ?q)Kx��´s�EٗLR7[��Vy���Z���:�gA�;%�L���k��0tDD]pᨏ�;����l�/����Z�ХV[�ϻ���t���MőW]��	 PK�����  �  PK  ў,J               113.vec��UQ���̳����������l�[�[�l��9.9,��9nD���S@!E�(AIJQ:F�,��^��T�"��L������zjR��ԡ.��o����ވ�4�)�hNZ���Z�mhK;�Ӂ�t�s�E��w�;=�I/zӇ�)��]} �`�0�aOcD����(F3���c<���1�n�>��Lc:3��,f�,�����1�,d�Y��T���+X�*V����c��m�ۨob3[��6����6��n���}�� 9�a�p�c�'9�i�p�s�����ey��\�:7��-n��w�]�q�<��y��S����%�x�����,>ȏ|�3_���-��=����'���۟H� PK��Uch  �  PK  ў,J               114.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK��4���y}�g��;)df���oi���N^��>�|�?��X�]~�3�����y�OϿ�����*��*3�����S�Ի�z��u.���!�_h*G�Rb�q�/�����tXV��u5��:��3���<u<����e�{'�}s�v������������׻�^�.�W�[UW��U$�aQ�.̼�ZBo��.SW� �<�/������;6�E�����I~���Ĵ�j�1�۽%�ՐU$��5�4�{���C't?����!�q��)/�zc��ү���{��O��3���	�3�j�r'����P���|��h�Rg�M*�WWw�1w���ʏ�-e��VN�-%��q��gz|�+��������X��D(��޻s�TqW�N�*�{����x�R��Po������ofOo��7�s����Uݎx�Ů"!�D]���E�u]�9s_�"�L����;�ݿ�����2�[�ͰP�.U>�7����5�3U�Y���!tOiLÒ9�ؾ�o�>y��m�������.�j�l�㪆��-^Ι�]f�+�E��x�F���?*�
�a���t��W��-�n��gw�qƶ���0Ӡ3�U���皷�]]v�p�(�ǉm�e�Ϲ'����㝛j��/�,��b��Ҽ3|���/x���3�3�\��J��J�++�$"���?���v���?}�K��-�緺X�MǓ���8E�iu���	 PK�/�<�  �  PK  ў,J               114.vec��VA���vwww�����ݍ�`��؊��
�`���]�G��s��e���O	
(I)JS&�G�,��^�
T���BU�����zMjQ�:ԥ�iཆv���4�)�hNZ�*�hm�FoK;�Ӂ�t�3]R^t�RtӻӃ���7}�K���n�>�B1�!e�SQ��
b�>�ьa,��&�\L���Oa*Ә�f2��)�9vs�y�gY�b���w,�[��`%�X�ֲ���86�m�7��-le���N�]r7{��>�s���0G8�1�s������<�Y�q�\��m�ȫ\�:7��-ns��+�q�<��y�Ӭ8����%�x����|�e�Q~�3_�ʷ(��\�����w#�PK{�l  �  PK  ў,J               115.i��UT���ni$�C:iq�F�N��������S���须����/��޻���k��;;����
�HQVA��
 �<��@���������������OF����OEBJHFK�����X�_s2 ���l�<� Qq>1.~��8A�����ç$ ��{|���,Om blI@&�k *1
1�S �|O����T4tL,l\�g�" *
*::����Y@'� y�+�I���#�t6���vr��cF~�\���T�L�,�l��B�"�o�?����+(�khji��Ꙛ�[XZY�89����{x��������������_PXT\YU]S[W����������?01�������_][���Bn�잜��_\^]�������?���E�̅������.T���c���$�R���H�����}tVE;��1�	t��Q`���?h�M��������o�y >�s�Ј`�IS�JX���;�����մ4�I�(O5�D��sG��@�Ҡ>�����־q�-�#�:F�8���C.-�U�����K!�%l��܆�z�W���s��5��@�
��0[�p��
�����ɯ��nk(��Aq�g~"+������v�ɡ�}��]&��9������IR�g����:0����[�@O�ːj|�ͤ�R�������4�Cٰ�o��H]y����d�ҚEHqa:E���2R�Oo�A3��rU�G�=9��^E,�w��d� ��� 9��M�ƕ�+��j�;��Vu4���//�7ifE�)go#.�:%��F���uh4M���/��q����+��EHZɢ#�X��LR��y�QS�ݼj���_�۵Y+���Yu�5F:��2SrC�}T%a-�)�A���<�N�V����G+��I��5W�U�������]���xYF8�\o���v���2R��.0T3<F�u�P�n� 
�)0A�w���i��n��'����_F�)�ON��P��<����� eߚW.���I�q����j���#
Nv����\S��J��u(^Zz�~)������r?ٟ+2�I ���ͤ�3�ܴ��r��0�͵+i�׭B���Ń�X��^�������k�A�r2�:�~�E��>XCV�k<��0Un��ŏ_�s`�5$����(�Q����#�t�1�gT=��r�i�&�@/��TX(ȁc�U��8a-�Š�Y�f����p0 ���6��6�~{(0w��;"���1^�R.�H:"���.ˍ�E�����?����{�-Z�ΰ��n�n\���~c��(�m��t*����sL�5���5�5���J�)���x�%��F�]�g�+�}�O���΁ɕ�����2�Dx���l:���Ә&]U~�������9��!?:Z���e��������ԑ�������R�bɺ�$%���l�ye5eL��)iKZ	Tzz���O� �b�L�7��N�Q�!�i����ڿ��2.��#t���@��R�(��jq��}%�q��.��i
y�fU߬,��	��'�W�k��E�("���"䭫�,���h��1"w5�K�LKb��h�3{ED(ˠ�C	|��&˳2�!]��M�/ЭL3�7��7�9��.{w�d�"���V����,W��N5XE���íw�p��۞2�S5-1O70�ZK��XŨKY�o������L��x�QrCE��3����5M�3���B�ĻX�����$�~��[����
d�ݴ����zX�733l>��4?lՃ���~���u\IA�W�~Ck���u������eU4z^�8�H��v/��B��T�Bg%�`8K�x,���VB|
�2���06̀��'����bl��Q����f��	 k�]f.�:-}[�^\
8���U�U�E'@xc��+��xj^�O�5ƚ�*��۾g�1�G��M����ә��f�/w
�w<[���}h'v>�t�^ћ��/�
S�#�5f$j�2�	#f��0�k�dׇ�yD���Mdo�zW��c%G/��S�o���w�ᢪ���@���L�\e�6?��p�}�F�����<l��
�x�k���eձ9;�e	��q�S9m��[>�H7������V�uE��>�)�aT�<�/*^6�̈:��l.f]����0m���m�T� "d�c�z<�����3«7R�"/;~W?�OW�~`�'��(�r]A��ߪ+���𥦍�� �2��.����E/��E~ϥ�J���m��� f92p��##O�t��
s\A�=L���p���I
�ҕ�1��Z�k7��ۑ�W�#|�oz�.�Yu`�f��בn�G.`��=�&�A��C�8l��O��&�3���0Ga������@J��w O�q�CKCh���N�l����2S���J1�o�)��5N2
�]}h�h|I{X�X���uC�,�]cg�!���P�Z6���yu׌��\���� �b�L>��P�UW(/s���*��q��7"��!�0���hq�g`�w�w�%÷' E�A)��i"MP��"��b�{ܚ�ǭ�AI�*B�;Q��ʍk����;_�]���ԨL�:�C�p'O�� *�/���#�v�.e��&��H&JiF��tX�hZ�����+f6|�UO�5O�������7n����&�'�Y�"��#�Ɏ����J��\��_�-�u�]�܀��Nk*}�67�р}Ft�3�8��B%�lsQ�шG��uCNj�Ae6�R�.��Z�ī�s������~�z��f(�o�(P��{9=_I$:�#�ӓP�?�)^ �qB�ƚC��|&��/J3��m�qN^k�~2�U}!�6���'�j�=�����{$͔��7�б�~��&ܗ��K����`JD��,3�Xsv�M����-=�hW%{*�e��]�����-/��+�>�{@��r���z��yU�,m����>��c�_��+fIl���_N���t��Qh��4Z�1G�	�B�$A�z%~�FjOG��s?�p��[�(����S�YL׈i�56;h&P����N�-�@�}������E������	o�}'���ec�.����wb�-Ձ�I�0S�7Z��.
�W}'�_����͡����V�e��(�o�N��I34t�	EeO��D���K^�����7�X�sA�����	�%����U��wBp��*������������O ��'6���/}�6e�1r��GΣX7�ګ���q�cA�e��%�Hf���u�Ɂ<�S��y,�Q��}�U�����o{���y./u7���5՝�Vg f�����!���L6u�}���E��������_���q_��!�jVs`h >����-��@#!�@���JٶSϸ�wV�3��塱\�&)�0��(fX.����}��z̘HY�}�
��f
��QM�q:��'z��@��IMd�^',�.����-��R���
��򃎋^�kZm��iL5+ۄ��\���J�"����{]�%�
IZ�P@W��8�r�ҡ-����B���SnU�̄�r�w� �PVy��������E�H/7�[�+wG�ﻎ�̌If_��юa�X	�f�|����f#!m\���yЗK�0��y��KJV��}�@^y��R��a1���*�Jv��`;"(	1L�u�qX������\07D���V�DѲh�sâ*x��?���^u���C=	�o���4]�#s�����Q"L�˾?��A?�P�.����@�b����Rh1���Z�����p���UO��o���I����N�8Ȁ>f=�/o�_͖\KI-3Ǒ�	t^�Gx$�<�@_N� '��]"ce��_�Δ'�y�
2}�J}��>\������^`�f�̚�f�K��J[���Y�hz	��]!KC�b���֬����t�>�]� ��$���6kj��=U�b\�����cu"������@s9��ʋ$t�v���upޛ���J/&&_�%�IGi���ϙ��������	���dϿP�UҘ�p[#&H[��s>��36u_��N�t�ü>8�\j�V��w�M6�x��ߒ���Iڛ�B�h����;����}�a�AP�3�8:�W��z��g�ܗHwUlqhs�X98.��_s碑3��C�"�_�S����*��:y����?$��;�r?��p���*�3��A�Gr�,\�"q�/J��]�v�W��f��d��/V��}�eR6Tqj���d�1�Zy-�s��l��<}�^<�ߧ��)�	8��.��C����3h�(>s���������r�sf����A�at�����B�W�vXg�%��tA���@�:R�@T[i6����Dӥ�"+o;��=�/��(��2Gi& H������ŭ#��Ș��բBG��nH�3O4�s�&,|�[*����y�G],o�2�:%���D�����>��&��a*vH�I�/PC�U�0�čҼ���q��N����L��8ʚ�`�J��~�ƢVz4�C��Nno�����)��5��/��<h�N�ok3q��`S�1�~�m����f�h�����Vg�؄s|��zLE�%1���"��e�����[)?tgy�Ͽfw�wÏ����n;솶�seZ����*��.65��Y�l lI��y��qe[�$��&�J���O�x��{��7�v�!�uh�@_�Z� ���\�:8�?O��^����n���j�t���B�ƣ���X�Z��$�^fH��Ó7��j�
@��2�/���5@R]��	��~�js�r�nD�����e���$��A�G�W�m��&c�{���ڐq����LR���!֞���t��G�����Ͼ����T�W�4�goP�rsC�M������;�^o�k�@8��7�pɸ�?��X�ݱ�y?�;��=Ʉ�q��O ������n���@2�c�ã�Ǭ7,�=�+������K��l`W��>ǡk�K���8H�v�d�X�s�Łܚ��#�Ōq�˹�92:��I7�]s*f��Ji��D��:����ސ��)D��5�շ�oJ��vt�I	��L�H��/`��;ϲ�y�y�1���#��d����U��(���k{�"�3s�����1�zW&���`��:[�>}�)��N"<���qe��!�Ҭ]▃ϞgM����;=,|����h�E�mk�Ĩ��b+J���aI����}�V����{v�l���_`��_y� �1�!�L��Rg�B�o�C��#���MM�U=�Ԑֽ��U��_K\�.��{UJ$>.�v4��Cu��������֒��r�B���J����� A�����4�S�t*e>�W�� j��3�ٙ��������*w8�!n��)%Mr� Tw��!sff�L@;d+x�፛m�*d��^���>7T%����Y�?���w�OGWy�9T*�I������-�#)I�����Vu�މȣXD�n	��_�M�.��ӨG�~r ar7�I�^+�qg�C[Eh�;���M�K�?	�z��[f~�F;�]��h���9�%�|\�\�>/Lo���q;Ј��$��EJ�:t�Tg'dڡeE��5��o������w���w��~`N-�v��1#�t*�I���'@��8���Ҥ��"| 	��	 Z���g�C@�M���9*n��-?�=� F�Ͽ So����+�e3���{���A��k�i-\�[ɿLIEǹ
�}�#�+]��К��w�a_�$��ح�ݴz�|��tAH����T�����|ۃ���~�6�<�&PU��Y6�p����x�T0R�?P��w��۷���K䀧��G)�F�� ؆us]�9����ሿ����ݍ��L��Bc�-���C�w��n�ݠ�pk⨜K�� t���Kv����Mx�YL�l�� ���ŧ���/J��-���dh��W���pW���%׊�w˷�����Z���Դ�����Ȁ�'@� W�B��I��:��ޫ�/�4,*P�d�j���q�bԵ���qQn��pݱ�kK#,��U����9�5þ��t�$��[�W�RBqv��M�e��?����G"�L|������ԛ^��h�G^��9w��`3��8r����닓v�Vڨ�G��K�C�p�����#eH�zRN��������4�e���&JJ1�j�z���3C���ѱ�F��S��Qڰ6"R��w��Y.u����mއ
X7����� ��)��jˋa��k��x$�E�|��57"g��R�a�V#���m�5~��@� թ��E�D��g�-֡�]�����ZYsF6c�1�B��|D��ߡ��\�6�<�#�������[����r��㢚���D��)�g����r�eF��)/6@;Z��&K~޼O���{�Ƿ�\��Cֻ>�f
~#�%0$*���	�CQ�i���
,i`Ġ/�މYƦ~U��u�X��� L�����,퇓nϪ��&�Pi+:E��U�D|�KQnx�Ut��������T^��Q�&Z��a���
n�*Y�����v�wV��)�F�V��"��.���k��hʷ��Q�f٬�F�����~��\�����CUʖ�k�2``v�V�@�;K��)���#$����>�m�KD���ٛσ�<�t�	N?�q'�3c}�A�}��Q��n ��pkK���떾�f� /s�2��\,�ec����F`M����)ђ��(.�";����H����� ���nz�9�gQ�泖��-J��������u9�W��D�ORq+\D�eĮ^�HfD*�q�y�g7��3)�N���e>�u��̠�ϗ�o&�l����>��a����)q>.�'܄>@��U�L �Y�cRz��$~�*�y|Sb����cH`�^�J}3��7l�[�}�є��kF��S��M����8��s��{�<6 gT:W��ɔ`�&�t}�U=�/_�isl���N�87����=�'U�^��/�o�F�
x�e��q����ɉ
Koՙ�{kz��PnL�5v�.w:�Bh3�`�����'��*�MJ��j�Uh�*�Yi���x�k�3�Q1�)����e^D�!�浸U~z�)�/�`�� ����{�����[�eYyt�E�s��g:��$J�#�xO2�K_�S�=�3��5�:�4y�iƗ[�����=(!�k�-k��a��q� ��bt��zFJU}�Ц�K\a�a��I0����V��j�D�/���T�pw��������#C�=���W�T��se"��Ak6{���/+�ڨL!�<����&�k;�m��U`zN�O u��t���mG��w��M0�{g{��m�	}%��/W�>"Y�=��^s�?}��.�;����	�օ�N�8P�7��T�1���&J����LZ+W�,�*���Ӯ���L�<Z���`D�5����ǐOd����S��I��!ɍ�z:���wF+`{_g�D2P^��0&�4r�֍B�Qh"���Vk��y���G���~���n!�ɒ߶�)����)r1J>���ND��F����6��(�/�KЂ����k���y��[�r�Ab8M��i.�VUH�\����&��s�`�?S�:n����ȴ��_��cf��,�����n��,��w:O �+�ҽ1���hX�Z6M����w1�������3�#���+���N�	L�)���m�v�'L"~�_�"E~���]�J�0k���$�K��
��:/���>��|Mٷ�!i E���C�3�sl|=��as�pfI���Q�ky�`:'�M���y�7f�!��1��@E�;���#`��Iq�/�F�2Ů�-�B9�˦c��@+{+��I��2`�"ֱ~1�Cc��'�.Ź=!���*�B��q1��Z[��e�_�K���4vy�ݍ
��@�Z�o�: j��h��Z\�bG꿧�|]c+B�������{�{)��6����=�J�6��_��1�(�u'P+����yֶwll�*ƕ�4L���Q�[Ǖ�º��S����֤X��-R6�\z/辥\�C��#;3J{�MSL�8Y���vS1;��=�cJg0o	k�@C�z1O��x�|�JvR���d7s$[�V��0�M/\	���{wy��B3� z�F]r%|5#��/�{8$���~��k�˒\/W�!#cO���{}aG��,q2�XQN���%�,!���!Z��u�?�?ة�q�TiԊ�L`3O�?��9�gYh�h�Թ˄k�o�z���C�ƴ�r��[���#�y�+ڒ�V�"�$ڍ������D�� �>��ו{�J��R)b���a۱x;�~�ډ�m���MW���y�{�q��}��3V�,�#L\N^(�c�����%~%�)>�x����#Mmj�>�|3�BS��B4
�����{��� ��Y��<ӻ�b�����n�']S���7,-��9���%�Cޗn��3	W1zq�
kGj&8O%�K��Mx��&P/yi�#��z7i��f��H��Q����~}؇��������v�đ��o��M�V�$�1af�~(~����I��;�1�$���_�%�l�tK��>�L^�I�<?�6�E��#E}0�&�1���?pDTz�NqC5_R{̢2x߮@������B?�|�}�%P����H�%&�e�0�3j�n�1���:�8��.�Z���jR�> =�-���)]����4�_PK����"  b#  PK  ў,J               116.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK��4���ys�m�4��8����7�d�Ύ4�z��'�3X���c��݁���T5n	׾�LcYF���K�H�+,˷`�ɾ��::>L�v��Zx���ڲ_{&��z��9߄�n��t��ٝ��~]j���/�qǾ�Θ�2.S%�g<g�IM�Pgz++�-Q0�RpQ���1=�3��Y�/���䥱h���H #��6��lեE-'��Y�����}ί��<��n��h�4p|�:�W�����EoE}�65p]��ܪY�u[ewZ��y�,?){�����&��0�4yZ�ɟc��g�}7�vP�c��H0â.|�y�G���f?��8���릧-n���e��/u�ڨ� �䟐pɒ��B�ֽ�(4oɗ@WV|� ��RO�$%܍gZ�{��9����'�0ԅ^�޾ڦ�Ӕ�f�/�X���㯫����&��&5J7�%��V�Y�X���;k����k���T�X�v-zx�p������͟R�ȟ�ucƻ�mb��\z�Jf���?��Z�)�X���#�Mڛ./n�'X}��(����4�9=��Ƹ-
��V(-�{~�s��K�w�t]�&�ʀg�ؕ2����4����	u�1_e�Ƕ�~]�0w�m�l��9>a�Wg�U��c�}�xC�ֶ
�:�g�:r��<��*��zv�;�+%������>�=�����U$�_a���P������<#��-�]�����g[�-ʤ{����,� PKm;_T�  �  PK  ў,J               116.vec��Q�3/����n}vwww7��-�b+�b+؂���\���63f"�,�_y�S@!%(I)J��(�E���Q�
T���B�T�<��^��Ԣ6u�K=꧈v�F4�	MiFsZ�2�he�ZoC[�ўt��S]���ލ���'��M�zo��0��(b ���2,�b��}$���2��L��h7I���2���`&��o��}.�����,Iy��n����d�Y�Z֥�Xo�A��&6���lc;;lv�]�f{��~p�C�G9�qNp2ˋS�4g8�9�s��\��㲼�U�q����}�;�.�����<���S����%�x������G>���E~�������ŏH�_�v�O�PKp�Jtm  �  PK  ў,J               117.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK��4�b�a�[7v�^��ܯ��暛�y���Iyg��6�q��o�[br�m�]�dʃ�,d��O-�����Kc��Ƣ.z�W��ϝa��[/����e�<o
��z�>Y�u���<����jO9nj�9K$�5P�U$�fw_�~�L����}Ǟ���%�W���~M����?�B�RZ2O;���	C��L��/��¦�v�ީ��<�m���B��ck���>�bh�/�z��iǿu�/����ںEeQ�V�=�pɭ3�=WΔ�����mq2���K;N�����z����C>l;�T��yLL����-��tO\{zJ��!�H�>,[�!x��f��լ��3����mδ�9�މ��� ʹSU���K�,�:]E��6΅e�s��-.��q���	��������Q���\�=N&�7F=^w#����,���vi,j:D =�έ��2s��2Q��_�1{z"O����e/�o�#�]��b���u��>����/l���kR!3�K�J��]k��o�"����v����^�<=���ҧ���6�`�s�\���<1�%���O<^\���x�2�������y��������n�9�3�]"�����1|^�-�Vzt�ḟ�V����6'�I}����W��sVPͬ \�]�����r[�>���[��$v�$��IW�E���Mw>|]��ǩœ����q}����ڏ�Ƶ��f.{�X/�lu`ss\I��}m�f���bQ��g�Ӽ��w��<#O�J����ek�ݵq�ל���8r��@��7PK<�]c�  �  PK  ў,J               117.vec���`����������݅�݅�`��؊��
�`������x8�qx7�"�$�_9��@qJP�RY>J'e����<�H%*S%+DU�UӫS��Ԣ6u�K�,��]�!�hL�Ҍ�p^K�Vzk�Жv���%���uѻҍ���'��M����ޟd��P�ei���d��X�1�	v�&铙�T�1��d��l9���c>X�"g�Xb�T_�rV��U�fk��Xg�^��F6��-le�mvȝ�b7{��>�s���0G8�1�s"��Iy�Ӝ�,�8�.&��$/s��\�:7��-���]�q�<��=���?�D>��y�K^�7��]�7��|���E�5�����=���O~��;�PK���j  �  PK  ў,J               118.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G)�EK��4�b�a�7�r�����SP�j��x&��{����.m�t���}{:?)Y�ݗ#����Rߙ~�2_EC<]E�7�Z�pBSk�Wkߢ�}�7�#�\~��|���M�j��Ɣs����M�`�r�x��<��zr#���8�����-!�<L�D��G}�٦:y���!3�x_	tUj�J|Ӄ�ެ�h-n�r�n���K}�����6�β5�u�*�E/�H{�#\X��c��^̶ܱ�*w���,�xNM��ub�o-	�7��u�+��y��U��Ι�OT��`��P��䥱h���H #�{�[����je}��_��4�'�m��^�oE�wx烈�WR�?�i�q��6_�^꺐]�T$���`�C��8�Z�)rZ�zÁ�'M�4Μ�*{�G�%�6��X�X��A�;{��!	��L;��t�Ƣ�$0��K��~�����A���1W��n�=�z�Z�{�^E&��NdZ�S��S{9�i�?�_MT)�z�����:������]�O��O�c�TWy2�r��#�w��ng1��S��_��{�z'�9*S,��`���㏖k��s��Zp��EC�����ً?�n	��䢓�"��?�m=_��y�Ӳmj�s��ͻ#ܘ�[kW��m������9V*�gO˽A�����o��i�Zuq��uO���]'g�����_�6��ƽ%���̥��������G~s�׼����+L�u�<U����K�j�,�(��1o��C��s��>��Tp�|e/��s��b�y�)��+ϻd-���۰����ڍ��ky}����Ƣ.\86*r�5�Y�_�����:y6-�o���Ǿ�<�*ۢt����� PK>���  &  PK  ў,J               118.vec��UA����������]��]`�؊�؊�`��^�{��e��+��r��4e(���\Q^�@E*Q�*T��S.j8��^��ԡ.��O����MhJ3�ӂ������ص��ўt���B������=�I/zӇ����݀�$���2��`d��(����2��L`"��l7%��T}ә�Lf1�9̵�'糀�,b1KXʲ��r��JV��5�e�ِ
��n���-^n���vv��]�f{��~p�C�G9�qNp�SYQ��g8�9�s��\ⲷ�"�r����&�������y�C��ݟ�4+�3��y�K^�7�����/�G���|�+ߢ�#ŏ|>~�_��O��o�PK���g  �  PK  ў,J               119.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G.�EK]EG1�0Kw�j���$����)�ϔ��4�%K��|RvuB\fX�x�ܻǈ�f��/p���W�"1�U�H�+=qnV����A�z��V�8[z�����3ܺ�|�����M�����b��Ga�V�QI.8�su�֎/*�lu�u�N��N�Z���m�����l*쟽4(����Ƣ��{�*g�m�>4��N��dm��Z������s�E�6+i&�t?S�ǝ0�Ԏκ��U���-��3?i��C�����W8�Us�Iٽ���w�=����뗳��<>�*^���`��jE�ui0���+�����ϙ�{��ΓO>�?�뺸��1�ݾ���V���"~�^����c��*|U��{�$�հU$Ё�5�Zϲk�$�Rv�J�?���3c~�zW�,��AH����G[&���v���*�E3	�1v�G��6ى
n�[y��uc��9�;-��>��;.�ԧ=^-�_Ʊ.��Q��N���.i�u.���2ui,��y�3��T�.�)o�t]�~���eMgGě0%�`��= {F�����Ibo.,���+�����Um_�YC�*��j��hW����#�VW�Sx�wm=3��fVv��λ/�]��{n���
__�՞t5�ly�WN���_�|�k^���ޔ�S�t�1T�-��u�徲Z���;7��7Y���;_`HE �̘�c���S���"�p}=OM���ei�'�
���ʫ���ŧ�k�����Rf^���&��<i3�z��Mёzޥ�<�D���K;��ky}�WO�X�Ņ/Px���k*OO��lhy��s����B��%���s��(�����& PK�|�%  "  PK  ў,J               119.vec�e��A��Y��������n���[��Vl�\�V��?��������DdY�?����)CYʥ�(oWA�H%*S��T�:5R.j���kS��Q��4�aJ�(+��z�Ҍ洠%�h�6�k���=�H':Ӆ�)�[�]�AOzћ>����d��b0C�0�3��)��F�c�8�3��Lb�����4�3���b6s�k3O�gY�b���e)��v+���b5kX�:ֳ!��F�M�f���mlg;��n���}�� 9�a�p�c�'9�N�3����E.q�押�5�s����6w��]y��<�!�<�1O���T>�9/x�+^󆷼�}>�G>�/|���)���!�ߑ�?��PKHJ�Uc  �  PK  ў,J               120.i��eT�������R�� ���0 (0Hw*5��t�НJ�t�� "1�����֍7�Žw�Wg��:�}�>go���(^*�)8� �s7���"@x�>��{�DD�Ĥ�HIHH�R�S33�3301�pr���31�H<�qK�J��	�����)	)݃t`V&V����v��8�@�K��G�s����y�������>!1�]@#�������w�>������S�{�*�p�Jǜ�͕��O�����F��_�`"b�Gt��\�<OxE��%$��_()�����Ӈ�6��-�YY��ڹ{xzy����14,<"2*1)9%5-=#���������������������`54<2=3;7��}qi�����z{g������������p <��i�G.�;.\||<|��p��z�'������
:�Tl� B��	��=D�"�i,ܾ�r��q��������������ZH�p��� G��{P���j�Y�=Q���m�h7���o���K7~��.�����-7����1�-$j��%��W�j�o�]�fh<�c���W-4(>Φ�Z�LKit�C�Y�%\�#K{�)5�\�v�dE����C�U�>��y���Ҹ�L��D��3R����k�ڷ�L��Y�	����l�9�q����$��tfL��i�9d̰6\�uU�ٞ����>c?շ�ߥr��˙���CC���W��RX��G�l�U�Ι�/,T��P�>ӀG��ʭ�Dj#�0W<��9��ٮ�څ��JV�:��RHW��w�U�N� ��ܸ��3˃	rE�]b�v�G��_&� �`�Y�GS�oe�Q�k�
���g���+�:°���]gg}�G�*��d�B����Z� y=W�X��7N�9�ݓ`
6��{�U�+cl�^�N�@+e䫷��R
�S���lr{{���l�Y��U��B�(=�e��-�nr+�R��Y�3D�x氆���'�Q`���y9 h%�c��[���&��r�I�^�h���'/�������u��kT�mU]S��(<p�O���3a�B��J �)%�����[ÂŐ��T��a!yoe��O��qA��e�'��И�D/3�SdA8��R��1�A�O0~�w<Y���ou���j�R�T�L�}�ʓk�N�W��O�)��q�_>��C�(�4��7�H�����XnM�ҋ~x��o���?sG<SfÖX��g�R՟���TU�)�����k�]��y�u�Mz;g�����_Φ^�y���Y�SXV���M�5J��H	�r�a���UI^$�^��%��~JO�3��͠���=�YWѢPz�q�]A9��w�5b�'�Ց�@t��wk�B���3�f�
�7<�?��2��	1�,�i��+�f�{�戼�
��d�w�Ύ�S�`��u�aԿyb��c>�o�k,�Hi�8 �ۀ^�lT�kq���3��7�����}�����`
B�V�����-@�|��+�!�l��h"!�"����0B�WaOT������7Q�i:��唵�mX\d���#��o��4kIl{.v��j����/lL�|+���#������]H ����mE��qVBb]�M�嬤�r`=g��vY�lH-�Fcz[�W;�-��z_�+�Y5H�i�+F�R+7Pc.��ސp����9|-qBP�59S%	������̩/8��b�	ʝ�j�W��)�:�0{�\X����Rg�T��L��4��K�6�G��l=kf�38�����l����'����-��5D�;gW��-eje�YO�ѧ�S����)k���P�$��U��i��+��e��X�:uD��(�P���ќ�����[YbG[m���� �Ȇ�]K��|Ks�U�*r�.�[���L�FC�_φ�M����Δ���d����[�Ӹ��:'��癊�č��5��3P��yp��	�?�.~(���泠��W�IW��v�=��������ͧ�C͌{�y����ȁ�˨	�oj��?Y¡�_�sn1��ZvC���1�����(ܤ�hO��������6�B���5%��w���F/�N�2�R�P(l��N��ws�AHW((Ib�/�%�8%#���;5����dtTk���_1����N���BǾ������W�7t"C�i��&�꙰��Qۮ�:����[nv�ÚD�Uk�}\$��͍���l��&���RFs���c�-���e��OW�a��~���IgE\�x'VM��ov�����w��9�tIV�s��[t�L	�"�I��fb��A?,����&��O��!B�%<�*0�NȽ��D#��0�j�J�b�GS�"����6��gU�N�ȴ����;�5���<���x �H�̡_,��~�T������a�u��.��9���L��,���%$)/�[����?pw�w�ls֌͖x�jZ�l���w�wn��Hx~ y���c�Vm��vT��QU�p3��j��a�82��
a�3zI�B��@3�3_��C0��}���Ü�TO�LFB�Ip�X�)=���2`x�7_�{��`�7&pPh��D>]�@���Q��Q*��4�_���%,�kZ��-��}����ן�u���LcK��z����@��������z�UH/t�
����%��験,INS9�4�כ�qSQd��+�6!�F�7���G��lǫ[ ��LD��!%?��������M|���P�{�Ȼ:c�B\���-�����$ڈg���-h������P\�ʅ�����B�$������ט����qy���+�va'��,%�2�Ǫ^9���G�٢���1-Ò P<M?�)"},�K�UO)������Y�q]�2v4���f�̫uZ�+p:����i��:��g�6j�2�{�WӾ�#�yЁ	��Ƌ�_��z7 �==u��%(��
��f�De��H�]iK���>ҽ���?�9k"��p�zE��U��gL����4��zo9K��n8�ӂ��J�ו�I}�~�P=]i2(��s�&��g��D�Δ3��N����I_�4җ��ʈ8���_�S�Ŋ ��7�2�Nq uJIi-�S����X)[�����,Æ�KɬA<d[��l�w��:����0#ٸ�՚{�u�q����za0+�#;t��e��<�O|K$4��<ӘU�嬶M��^�����I"��9�m"�7��&�������9)�yÛ�g�,21��S��ƅ_~�읗
+|��u��g����mg��3ogz+���uHʇ��P'^�B���v�����{�p�@�6�,3_�қ�ᗆ��3^�=�|n.�sJ̇��!���:����/Q�<��æ�-1����^T�%�ؿ�TH���&[��2,�ϱ/n�=X�lAS��Y�Δ��GŪ�v�O��H�kl�}ğ��]�˒hV� ^꼸��Y��J���?����j8��(��S������÷@��ߪ����������N!Y��#�,�PM�R��ɒ�7�0�'�g'�=�l�OQ��qK�Z���a�f�&��f�Ӓa�ˇN�&~}G�^7��&/�������*�Z��<�O��c��	�V���f긽(�&��ͫ�z��06%�mߢ+m�#K�+����B����V�R��<�z/r�z[e}�h������Ǹ�)s@�H�`�їY��m񃀮��=f�8�W������z)�*M9Wv����P����2�-_4�~We����P��AG�EF�}�K�!P	ߣ#|2�i��Շ#�M�_��������~M���H�6�'���.:�;!��l�e��XիdHR��r$^�V)N�CĸA�6_Y���?��^~���P(H�iPį5���\�I�R��k\�'�3�b!�{0�#([)w�2�3)Uy�j웁s�R�~5�h��pLmW��cq�-�ٓk�3嚋������%�p�	���oʿ�_�SN]��X����or�s��p"@h�F����M�ո�ܡ����:=�_��ܐS;���È|���٣�hTjh~�H�	���ݯ�X��`p�QB�aY{ Fڠ$�%��L}Pkѝ���*�z�qX�;�:ѐ��x^�ӝ��j�{Ey|PĪ�OE�'��)4Z�[wb���G�hA�$�弲I�\^	q7�@�v#�B$�T���[(_ͨ�fo�	k�ԩ�=`s����zUlО=���3��BQWu�m��"�/�+�u�Fq�T�4R{[q�p$���O*)a��TM9�&>���ɧo���]�m�Eɨ:̀��Q����|��:vy ㊡��آ.p��h���\9��#����l�~�W<jr�Hxe�sI�qd���D"܉R�쑅;v$
U/�5�qhp.*���B`�[�݀��C��R���@�;����kU�p�||�3DP��h��M*Z��w�͐�[���}3}E*nvH��
�����`���d:�{��t�o���V�b<;�NH�/ ʫ0<�t�x1`<�eֿ�"*|׿�^wS�Lb���͌�R�ӳ�9�_����AS��*�(�⃺E^'����Ӑ)�!W:�i���T�O�JT�GZ0�ȢX�8�G����]Z����k��T�-�����d���n�`k
�Bɛ�rQ�[��:oW:(��� ���b���~��;�?K=���-����pSH)t��<P<dS���ܵg4��.9Z�C�8�ꍻ�]�MS��(���e�&I�z�5�-�r���+�z9���#����6�U9��(�F4ɷ�߾���g	�L�z��x5;n��:�3Z+WG���/h���u�{T!rNŢ����F�ɽ��}5��n���9���`*E?��yk�{�5�1���婰2�so�UE[���3�Rv|J���I��c�x9�%���4:��P�\�w�g�?���
뿻���Jp\�K2�52/�ʅئGU񣝤�.Xv0]�S'{݅��O�����FZ����b�k�f�֎� 'U�$�F�E/�fy;-�|x�W4�Ѩ-{�� #�z~�%ނYA��i�,'9h�~���8GT����M�e�b�yxB��Ȇ0��.ѪN#=>���x���z�p��/hMgY*�/u��},�HoW8n�ǋ��T6�Ñn���Wh�Al�9ͳx7t��<��K�و,D��񛿄�H�{)�_��x����3]LL��vV��º|!d	L�Z+�sJ�&� �F���8�_�<����7d�	�3Ky� W�`G�_��:L����Vd��^s����5D\��#z���&�w�ƞ�iA�J%��mM��5�e��!,z��[m<b���Wiak�8���_�������k0��
�V�ȡgN�����>�)��{�<�1���&U������$��'�-K�g�n���ށf��%d�֮�;�%h�N�xB�����~yd��+v��;3x��E�`lr��Pj��!<!�_>�l����Q�b�[x�6*���U'8�Ώ�g'�,�e϶%�\_�u�j�-y����E]�����z�3`��lp�ԃP~ǐl��'YzNn�lb(u����g"ƴ��J]���W)~�X�%�$��0��`ł����
ȿ�,5�����e幽��������\͛J:ز*�Lm5, (�'d/I���	�8�������t���50w��� F>�D]���s��E������/\͏���KA؊�8R{�ԉ�~����H���ύ����/\���,�0�����lalP��M�a����_�ӈ�L���µ�R]��t��O
�M�[�S�	��=���rj���iS2iVH����,q}�^&6�Mұf�Py<^D_��]��2� >p�]�_>�r� ��21A����/�m)��(gs�B��ґ,�w�t�#��"��t�(��x���~�M5�Pe�U����e�zÐ*�����j��v��~s]5�@D �ܜ�/�%7���M5�ߦ��=��}�M�;�㏵�O�j��~��9�`te~,��K��i� ����֤�� �3���PT�E)vC��fܘ��&xM��a���A�B@���W�Ge�o�ѱ�Iz���+$�8[��%1{����$w��@�Π��m{>O�*����2�L�&[�?�3@�T� ���1z�.-~
�4V����&Z����Sm<\��2�:: ���l�G��ڧ�ߗR!��������(������O)H��{��
_���"`2CHw'��C�&�WxzPS��_�S�<�0^������
d<�ɥCr���ȥ�ubQ8���uũt7�p3��Y ��	�R��*Tυ���O؊?��P;˟%�Ƨx�o�,P)vo�Rsf��Se�[� N���~��hNQ��v�[,ڵ%�����hv�Sf��+�ةC����@<f�f��Z�2���Ж�y�Wi�)�U��j���Q�b�?��藽�~�M���~W��Q�3�ʥ_+}9Y���Z��"���\?�� ��~4���=	�4�����>���;j6�kI?��	OE����qi6[_�e"jBtw	�q!�=nxH��G�y�{���)_!�I?K?%^���3���*y�f1�o���&�ȡ��=!��ezZ��{1�L����|��a��������j+�Ʉ�U�N��\����M�b�/o	_�kZ�����Ήk�@��ŀB� H�X�������ً�!,s��_ +���y?��{�_�p�*~4j%S�ʑ!��xb���[A�ۇ�K)��ѩZ���}y^��Iz��2XΪ�#I��J+-6�_x��Kc��r��+g=��E�uZj�w���в���N*��0_��f�+�7���ӛA�yF������:�z�LSUr����,O�JS�z�׉+nth��p�a*��'����v�X�` �d��2ϰ�4l�*�"�k���1�6���h����ZU�E�2Pm����#c�Mې��3�t��2�A�q7b�\w�ϑ5yY���M�^[�g��c�gwh��=*۸L�o})���Љ1��抚�R.aR~2�'�fй�I@~, f�~e򏹇\i\r 7n�e�x�O�����SN�[ .n��[��X���Q�:��?�&}j9ƭ[�p�1��U 3��C�b=#F�R|/Lr+�t:9�),2�S��H��}�X�do��t^��E9+�3��|N�u�8^Y^4�o��T[������klX�]��eUQq1_$`C��s�@����5R�Ý���i�=RM�DW��������&�J�u�����A1���J��.=���V����o�+����2d�M�{~8�~����&���^P��)�V�H��ء<r�njD���v'��q�VP�ݮ5�Ԯ�C|��<^4�$1i������W���a���~�~�GƵA��_�)k�t��E�tT��/U��������cq��"@���[�J��-�`"B��f�3��3:C.�7�C��ߠm�1�v������[Lg����h��ܐ��ox���.��8g�$�t�����5;�B�H�Lf��c�o�_��ދ���b-ϫ�S�Y��<8c�vZNW�|[Z[�i�D@>��m-�H�����X,dOL��K�,����i~ ����]g�wy��}?�����Q��૥�;π��x��.~�	3CK��/5:�GW:��U��U���Dv��W���
|l�:�#�F�V]�L�W��Ҵ��8��O	�!k�3#H��I�g~�P,���V������*\���� �*/z�̺B-�C�2�T[m3-Vie'��Hɰ�~�"�e~f��f��/���G���1wT>W�k��TF?4�i|�2��Qp<P/�p�f��It���Ց����T�8�z!���m�c}�S�L��z���O�K���1���HW+���.��g6L��
_D��K�O֏+<���}IX�u��$�9/��:4�=�&[��sn��̽6��&�RMa�}�R.�>l���ܪ{�� еb)b�/Xi���3W}{��G�9�H�pPD���O�V�����cYo�kF"����%G	���muqW�4Y;��Xt�m�;��/x�'U�Q�泉Wń�L��+g��mM�^�kY-�w�����9��|�[�rNo[NB�ky��9�����\��|wF#XWd�K�=`����(+��,���N��o+����^'�v���H�<GP��|R/*������q�yz-���'��2+���y�j��z�s�GB%L�l�T�KF��뜉^���@*��x�w�ΊZp�11m!���XKK�A�j02[k�j*({0H��t�~�z��ⁱ��K�����}3���ɝ�	Pn�N��pc�Չ;��4R��{2�F�Q���4�/�b7Y�S�E�C���XK�BLEb,<[`�U�4M�q �;�j��%��.��ޕ'+��ie�s�(u�g���P���S��c����D�,c�nK�4����˷ ﯴc�3�����)�37U�
�h2?+X��ܢ[�K��xYZ�|���S�۔�Ѥ�@/鄼���D2v��� X1'u�?<�Q�̂�g=q��Qb�t3��dV�O#1��?�%~-��jY�r�k��4XD��B�k5_n+j��ЎR*#���e��g����FM�㏩����d���%����Wjk���b�Tjs�"j�����觪V����[�Qs1wmZ�Q�).��WR]\�O.r�4q)���Zd�(��=�ڛ���	���
`f|��Y;���@Al���,i:���D�Q0�����PK>�M�"  $#  PK  ў,J               121.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G.�EK]EG1�0kG��풢%WO�:-ɈsStj���hӬ7��l�X��o�����aM�$�N�����	����OMm<���Ƣ�"����Um/�w��߼���Ř�e�gR�ܽC�ߪ'�<u[���imx-��0����f�	��cL��K��b/̨�PeU�"��O�B����nQ�dd�<orYQ�H��#� c\S9k�B� �c��g�o���q����'�抙~������1���kS�m��>e��q�B�ŎS��ם��S7u{q�Ǔy���&�:����������/L��X-�*3^��m׾+�[$د�n���������,��x̳���ɓ*�RG�,�1�˚�^0�Kc���.<�y��}w�<*s��^��}C}ԓ��On_�v�g�2�����ĽU�}kg=9q���g�Oܒ+��FM]��`��G�����*$5����E;~O�&1�J޺�8qn��zWO�Y(��_������b_]�Y����X4q�� ��uw�Z��3�0��`hg���c�{�D�FitQ�{�[����������m�����s{|vx"w\���//�,g�`��?��� <`j�Cj�L�㮎��@+���2��=w�V$��R�a޾ܱ��hS��e�=�˚��{��O�3
]�u�6%�y�˝sjL�R��i8y�$n���{���ul�X�9������+f�P�6�����7$~}�+|V�T��"�w��j�m���#����N��[;�D('�m�N��e�[�-�/�r�r���G�C�/���,����^�-������z����c����m3��嵰��MF�nv{\�}������45�m�ߤ��ba�rf��ͺ�f_�O��i�e�X�*��& PKz�&�/  E  PK  ў,J               121.vec��a�g���n��n���.��.�[l�V�t-��?���G�ý0��af"�,����e)Gy*�¨hWI�L�R��Ԡ&�R.j����R��4���4�qJ�Į�ތ洠%�hMں^;��z:҉�t�+��"zd��������/��� ��YA�3��c8#ɨ��Ѯ7F�8�3��Lb2SRS��ә�Lf1�9�e��|���,b1KX�2�����n���լa-�X�6z�Mv��-le���Nv��=�e�9�Aq�#��9�INq�=�ȳ��<��%.sŷ�*�q������]������ǔ���<����%�x���.�������,�ğ�)�9�]��'�"�#�PK,�<d  �  PK  ў,J               122.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G.�EK]EG1�0����Z�g]ڼq��..�6ZM��j����g����{,������O<�9��l��Z5���`����7ں4����lO٬:�'�(�Wf��)�N�>��q���7l�S��_��;�yף�5�ss/՟�\�3��:��N�*�����������xēYҚ�끞�O�r{���Ί::�q {�ӃW�l�񩹣iy�t���3�T�זݺz�*I#�cN�<r����jX߶۲�=w�I��N�Z��BO�1^a����������K箓�ix01����Y]�]Ep`�k��a�^�~<�K���IG�clf~�-��#�l��S�1�O��\��tY~R�n�|�vW�`	<&�M����\t����#����Ln;Z�e�)}a֫?��:��|v�h�q�> {z���7W���:uY !����}Z|2��X��w]�,);*��z����S���W�:o����uC��E��SM7GO_��˭�PRض���k�\�֐�~�C;��>�:��g�P�f�9�X�t��_[��tw.뒜D��L��7~k0lb����h�����=�omd�ylc��nk�6_�����nr��=5Y�KcA">7�w&L�V�:�T0s��O�V3?9y�Ջ��b�k�KU��g�=ΐ��s�Y7:�U��h��"!�8��`'wk����+LrW�?�_}����G������)Rޠ�w�q�������ޅ33LrX�_�_t�J񹋵�N�9fg�a��krض�%�g�}z h_Κ��	�^'W)��NV����^`Xʜ������}�ع?�w�d�,�N�U��cLR��^��e]K�F����Q{*�7��q-�uXޒ�|���g��?��kQ��� PK�Jt�  C  PK  ў,J               122.vec��Q�w���n��n���.��l�[�[�5�l�ԧ\΁{.�DdY��P@!9�R��TH�QѮ�^�*T�թAMj�\Զ��ץ�i@iD㔢�]S��iAKZњ6���vY.���H':Ӆ�t�{��a�S�E1��C_�џv���P�1��dT��h�1�X�1�	Ld�����j7M��f2���a.�l��,d�Y�R��<��v+�U�fkY�z6P�n�6���V����d���^�����9�Q�q���TV���r��\�"���^�W��unp�[���]y��<�!�x�{"�R�3�󂗼r�Z��-���x/?�O�?�/�'�F�oο���W��w�PK�ǉtd  �  PK  ў,J               123.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G.�EK]EG1�0���~I�>�������~+.���z�KU�>�����E=���(����i�+�IN���x��DE������4��/\K�7z�������s����e`�"�rk��ʙ<��1�o�3H=�{�p_y�Lʼ��Q3z�e,�Z�*�Ko�(�r��lǉ�������͚�����ٝM�����v{x���s��nx{m��[@|_�϶�ڟ��;����\����s����L�ξ�s�4O�=T��c���/]"5ŀ�H��\�jn����z��=3�7$0O;g��cB�ۯ�kNݚY�)x�D�s��9��O���w��R�O�үZʰ�O���:\��~K�\�Ĩ�������O�'ķ�9�p��E]ZGD]p�R����҂e�����y��
�Y���V�~^��g���'2}���%g�[ֺa�G�����
�%��/?�z�I�B����������l�}7���=�Es��m+u��4��-6b�v�?C����iޮ"��Rƫ�����R��<uQ��V�1��y'*��+ߑЛV&آ�׬��3Rb��SM7κ��U$�_l�����1[�=۵L�"�W{f�����*��[��[�[�uhO	y'��y�V�.�s��V�l��HX.��d���݅�ng�w�9<��/�lV���O�K���_V5�������O���S�⭛桤�H���������W����Q�U|v��1����ؿ�a�6�Fǻ���<��U�9�{_��}�k+�-T�4���ӖǗ���w�*^�71���x�t������g�--��i��+�ά.�ui0��L�;E�;�46	6�ڨ�c�����Rok��<�H[oEK��p�sB賌���DO=Ho�����K��W�
�Kj��vJ(�r�W�_�b&�w�U�_���~m�����?�
^��I�z�t\e�ɯ��T��� PKy=u!r  �  PK  ў,J               123.vec�e�UQ����kwww���ݍݍ�`�؊�86؂-����l�<�g����e��QL�<e(K9ʧ\T���W�2U�J5�S��)��j�u�K=�Ӏ�4�qJ�Į�ތ洠%�hMں�]�^�@G:љ.t��SD�,%zOzћ>����݁YQ�3��c8#ɨT��Y>��c�x&0�ILfJ�b��4}:3��,f3��̳�/��E,f	KY���7Vح�W��5�e���F�Mr3[��6�����b7{��>�s���0G8�1�s���ʊ�<�Y�q�\����+�*׸�nr��ܱ)�w��}�G<�	OyV��|�K^�7��]���>��|�?�5R|�����O~E!~G�PK��b  �  PK  ў,J               124.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G.�EK��4Psߚ��M�ǭiQ5�#�E�>�g���n)��&{Gۂ�WZ�"ߢ.�@W�QǌIwʺ~_y�5WGlڶ�_�$0�O���sB�_�){=�����g�'j�LޙG�ha^�,��?"�3���)ڭ���u��b�2��=�����r̾�[���fVui�R�X�ŀ����2;b�������?�����:�=��[�
댯
��ݯ��鰬J�;�?C�ه��9Oxzԕ>�����>�q�.o�<��<1��'�\'��q�D��󏋸N��r%�� ��pa��YW��΍��3�f��ο�1.���Ծ�vm��X��3=k&��������
?o��xc�����+�]X������=O7�_ﺸc��k�ғ�'p5�S�-���*�����/)uJ�ƭ�?��fR��=�|~�l{e�޲�6�S�	{����N����`���^[~]�b��r�+w�af���K;�J��-�S�6�ރ��KE7ݭ<�o�ӟn��<�0���줋�""@G3��%ujW��5�խg�WmǺ��?]�����[*�"�o�|��ʖ��s<�S�����K���!Bi�^(�Nd��I���?��ܯ������,�Ź��z��p=�~/�6����V���3�N]�+zGB����k��ٗZ��"��q�ꩩ[ؕ�ZK������ڞ�,F��bE��5)Tpub�P�`�s�C��B7?�>��Z��${ݻ��/7�
�|��Snk�yV<gܞ"���D�Յ�g��|��Wo��=Od��u���.N���v��_����>��d�y��]��R]eVȯ�;ہi! _��?rXNe_��S��
���:kx�ݞow�gܾ}uSq�V������q)�W�oP�{����ʵ�e����,�fz[gNC���K/���dᆛ�l�� X�2�����M���+�y��t�Օ�Ņ�ҽNZ-��o PK{���  �  PK  ў,J               124.vec���Q��=g�������V�nl[��Vl�V�[��S3���bo8��e���P�y�R��TH��hWI�L�R��Ԡ&�lj�:ԥ�i@C�8�hb�ToFsZВV��mS>�e)���H':Ӆ�t�{��墧ދ���/��� ������2��`$��
1&��X}��D&1�)LMYL����`&����2��6�B��%,e�Y����n���5�e���F6�l�[��6�����b7{��>�s���0G8�1�s����tVg�Y�q�\������Uy����&����fŸ'��<�1Ox�3���K��׼�-�xχB!>�O|�_���)~�����͟(��H� PK���D^  �  PK  ў,J               125.i��g4���G%�ed�N��ѢEg��(ѣw�K$����QF�c�Q�ѣ3^�w���~����q�u�������0�� y����� 0�P ���@<\\\||<B���O�Ґ�S�ӂ��ӂ@,|�L<� �'����0�]BF\P�OHX�?�`���>!�~��Z��(��� R<���|,& &))�C �X'��&6����& &&66�c6�1�&�!c��k[�2�S���1���P�L�Y{��P=���eec�����Tx������ZWO����jckg�����󃗷���xDdTtLl\jZz���/_�
��KJ��+*���[Z���������g�ȹ������[�;v�NN���_\^]������?���E�ȅ������.L��\ ��a ��i�Z��3	��Qȧ���3�SZ{LP������������������Zba<� _ێ;�-齻SnE���,��W��I���b��f�b�m��9�[��`��?B��J�L� �mMlg|��F�����,O+�|nN@�?V���KQc3&���3MI4�WGM�(�CN���r�2a�Y�����SOj�=-�c������/ 7 c^�����ᗒ£\�8�o��I�3[�Wl󣐸��ҽ޹�Qњ�ލe��a`�������X��QV�����6�k�K�Y:���n��>��'�s;��9d#YKb��Y�4jy����[_��v"WZ�j\�9կWj�/⭛�P�S�Q
C)����3m�(��B�=+�.�ݏ@���,� }i�#dU?�����j�l�e0W[��ބ6S*����Ye��e=���!��W���C}1��Cb��P���t�c�:�����ں=9�y�R� �����Γ3Q��b���T�rjp���$wyi��_�|�$�>���ۀ�YQpv�ZR$����},�ɂ&Q뚨T�.�����ƶ_��7ESN�;�O'�\��Ω?B�p{����&i������f�3�N�8�4L�z�\�J�/�̎�D�&8���Y<���a�Ѐ�<�g���|�Ϧ�u�ώG�Q*������T�K���^�t�mc�{J�р��Jc��@2fÞ�j��3*�";n���O��ҟ�(c�]�_�'���&;�a��"Ue��6��;V���ru]n���$�Ρ�;�v|�������o:.�u-6�p�1!r�
k���d�'�+�cYf�:��J
�}���'�`/=�EvǶ����N�4v���C�9�u�"���'�f��y�3l��1ω[���UP~�y7!�>8�Wr;۶�Â�{�7�e�������E���ʆAߜo;��Z�M:��_�p����!7?6|f��Q���\�X�il�q��R���ܗ���u�ʋ�7\iw�y0���b۔6���6i�-�PJ�Q�M&��`^n�_�����mՍ�@r�8�t�QHh�Q0>��5�QpAM%�N��vr�nN̪��t�в�p_!#3�q;�qR1���
�1I����5�C���<�RфD���T,��=�\�@���������Yۺx��V�d��|�����2�\���EN�2��>��I�@D�Q]���W�ȭ*�4�@а��&�����X�'N�~v�]�,�����E�S3L���lS�朗�k�����d�u��GsK���ju� ˚��*c�4�n�&�4rU��+�!sf&���xa)�vhݶ�����c�[���*m;c�Y�+5�Yʲ}>y�I!JO?�^���T��#E�E�����٧f�_���q
�|=
8�y���`���+�x��2qV9��H^��CI�"�\�l��tH]��y�v�+�u~�>�?�Ix��
������T�E9v�eH-P��dy�E�\��lcm{�؎�!;��»�[���yם�]���MKH�6���	�y�W�@���L{9��A7V.D�q�R�aZJ��_����?�fsy�
Tji��8������? � v���]ݯ��^D�||��l�k� ��≔�����(i:��~۞69ι[�HX{��Q�������)hg�3s�?Լ^	ȇQKof�])]J�Ґ��&U���R㢱���.�^�$�-8gk�⎊V7:Ӽ���
�L�e�t��ӫV�շe�����i��ה.6���s�"�f����0=��Ҋ���s.=���(A����g��z�|oL9��0ѕ��r��+$�h¤H���ȁ |��Iˀ�=o�g�I<Z�(�r1�d@���H�(7�`��n7�)&�1�F���4��W��@x$z�[�(�[�yDȮ\�dϺ�Ip��ώ�3�����u��@������7����<� �a]��_]o�� _i��F�$�|^Y�}9�0*�������d�o�2'?��_�c!�:E�>q�TW\@Ni�P9��~����N�c]R,w%���_*#(.Z �C����6����,�?[�^b��͹�Y�2��E 8X7��%���a��DϤM'��	E��m�AC��Q�[J�^ګ'��7�F]#sȬO�[VvH��.Tu�$Vx���p2Ԍ=v4o�ĮǊ,��n��y� Yy ���į':�-
�rs7,Lt!��?�7�w41��5N���� ��9����S���(*�5��"m9���IL�^���g3�]����L=+��{�gjI~�A1��H�8�Z���H��J�f����d�JZ�Fʖ|p����_7\x�}�m��W#���J�c�mN�L�l-y���Ì�9v�~lz�[5?�>�w�i�*>..��zu�m0c�Bf>����8KF7�xb��j�r�Ş��;���ۑ�>��"�����G�b�3�h?��d�C|C�״�r��\�=�b��~ 4�U�W�@�mU�O��ˬ�ヹP'-���)Ú��4������[�k�@��ϕ� ��Bg�]E��G��i��o}ӺD]#DaaJ۰�Om2DHpre@�:Ga3MU�_�����[Ќ�7�#o��)�7��q�!J�2�&�J��͓
�T��[����I��F�'��O�������U�_�d��d��V`r�鐳�[��:\nSw�j��wlYdKܵ^+��1
��~u+��CCjp��S��V`��2��1��P��'(�֯sYȁ ]A0�b")��w���IG���d���S�}�O��	��|,��E�_Mi�+w�L��eLTF��x��N�Ի#n=#�FK$�C�;�MD��t�������p��������)�����/4�������Ӛ��03��E@i%���7�H���t^�-�'�#  ���?�$��������:�iKӺKVc��H!M��Z:oq��5�W�c �`?e���/�耖i�������C�ϩ�	%H��:T�L=���Q��X&N&n.���7��<����:�>����GX��_�4�Ք�i�{���1O��4q�@�5%�r�j��^F���X,��],�4�V��=��
p6��k\BqBzp�}(jKU�U�N���7$. ��]�>���u�@����R0o���ި�N���@�t��")�j<P�@;�i�f����;���U�Weπ
<�)�&�.���ʉ$�+�z*�OR���u?-��!�-�}��㿶� �o}S���E]V���3��t�yY�Bf����R��ס�N��s췿�5��m��<l,�s� \��~q�y�v^Ŕ��Og�?b�<s�lX���$��A;���@�Y�j�]X���&x�4j�Ũ���O����񯝄�o�{�}�7��b�	�R�X�{ ��%�H��Hp�|�Y� ���Ǎv`M��0�xlFQɰU'�d�	������������@��3(�W#�4||�@%�k�d1�~(>4�|��$Y��4���y]���(������������蝹�m���>���:_�D��0����Ǯk/VA������N�a��? nnh�ռX&�r�}~�MW����h}={����^�0���?Ջ�ZY)b.��IXe�s�(񒛱��>a��b@���:,�RUSY��/�	��J����9��<�oPZ;�'O�g)�L֭SSm��HO������.�;�19�5��B�F�d�> �Q�O���	����D"��lƗ_{��X�'����Oxu����NF��
}��kZ�0�'R8���Psiʴ2���˸�o}Y\����	�O�zH���,��X8�0��|>�����'��!:��L�~�mi�D�X`�;����U�O�|��-]ԣv�[����	Mz����Ƞ�"�R�?�l��W�TiicYJ��+�U�D��s�O�(�V(h�:�Gfk2J�;�����J��,y<.o���\2I�.�����Y���=�fU|4���d�50u�\���$�t��t�~�U�6�*ƛf�v���W]��#-�J��҂���U��2G�w����Rm�W]�^�߆t��q����-�
v1�oxR��nGzm�Q׆Lф��[5��lՇ.��� �E��c����J�%����l��Gc�e����������42Vx����YKmnn7�i�yeŰ�N�p%
�۹�A���S.Żm�N�@�#��J�Sw�(���\	ܤ�]��k�ם@�>���鳛G�[��1�r��D5\��Tr�pb�6��o�7��Ǖ�w�ė�Z�Z%�>tZ��XQ˝&�LPs̈?�Z돳�ڐ���_�H �>�m����~�aRw�=wq�z4�#YrgW������uK-��60�5Yl]��X���j�����4YA;�'R�rʯ����RԨ�rk�e����x�"�1�P(������Z�cr3�|���*��Yc�,&^�ߙIP�\�Ί��6���_
�?���x�B+< j�������Z�w����4��UH���
yTR��d�Ş�l�됭л��y�}D��%��	b���m�k�}�p�r����&���(1i�GNMb:�`�MN!���"17/փ�M��~��@���PuC̓�=.��9fMyk��b�%�ZqO�#d�Z'�	���&����>c���6%���,���A��g�@�\�b ���}T�����3(E	�I��[i�"�#�UJ�+���L�{h%�F}�1&D�/�
�nz�j��g�Dk��	u��
��8���o+�-�n۠ ��Z#_G�e�� 0�Vu%�bOH�k���E}��D��d�[��5���c&x(�(��_uO����M����:��)iC5"H�ɬ�v|Y};�\��� t�=�ꏳao~s�05�UZz�z$�y��$.d�r����]O>��|i�{�ӽi.ɼR"��Y�(�.������Ы������IpE���0G�WK"���$�����52q9s<1�ڈ��*�u�o�@��\���O�W)���s��c���L������2g����K���� �K�Y���߬�_g/�C��UT��=�:��-t��u�P�.~�2=������3��{O�eǴ���d��]��Fk%5� �]�W�c�6zx:
T�`�����3�
'����d���lT?x�����ݸ����(q�	p����d��İ{����t�k��){�ͳ���h��U�ճ��|~�#d���g	on��~��K\>�ŵ�z���Z�kcq���E�׍ M��I8��ϔC,���F��5�J2��.��K��|�z��v/��Ćz}r�w"u�n���aS��[����2 ��DTY�W%�3��q2��(>�#�~�����c�'����ƍ����%P���� �J�)��9��������(��%�r�d\]��Ȧ
���RkA�C�|�+* �r�'jB�y�_0� �Q��IW�M�=�D��T�.1N4i�$�H^RuaV��r�T�jǝ�#l��^��m���JT��T�m��fu)��*��w�h*<���������#YF���t�6W�RD�$����{�؄��w����� �m'Su���Ӕ%��D\�?�m&ʹ�S1Ǵ���q��76��tv��9�egу��dԳLW;ic��2[q��QL�$FM/i��烅�&
�Ae0E`�T?�>P;�M�=�)OW`������
?�������uS������9����%�f���]2(� ���ߏ��w�[�k<��}�.F%�-��ه�wj����&H�<C��LD��u��C�VAz�Ub��3�Jj�[�2n��q�c?K�6'�y&"��eTǄB��sH��%cں�'u;�����5���s3GRO��@v�g���k���?�{�ā�F���	�X�ߩ��'ˣE�.̷V�
ӕ�����y���7N�<�{�&%�����^<���L�L���a�(���gg4�&��!�����Y|��w���ߘ"Fߟ@jڒ������+��d	?s��q._��]�|x�/���%��u޻^�~ο=DD���1���aL�\vI�[�����Ҏ����c���S����Fg��H{"n����m�p�I�,���*��F���i@������kd��д�Ey�ڤ|�a�?�����Kꃦ\z鳉��~%2!|��ӥRYj6��	�-3���8��?���#�4���
�<��6w7�5Ԫ�({2�����۪H���&)u����\�3 pH��2�=�4�ͳ!�R�Ax��3k~&8��6ɩ}ngD����Ch��F>�%��L�IMdՏl3��6�Y���"��4@��]0��e�x�?er�?/�6����:"�1&&����4C�o4�)q�D`dti�7*?��&�oDN���g��8=��|���8���di�����~�7`Fe��<��A��;��eq�Tc"�N��0�a!dI�����	ءhE���vL; ��D���$i��H��E(��f���+���̹�����b
�/#��%�+҅�;��`�ӷ9x��>����w"�+f�=����n��M��#����<�}(�ۖ����=)o��Z>�=����՞���)����,���%41'�^KX�L5_���_I	��x�O݊~���,t�]W���?��|qm��@IȩLO�y�)��*uo�JY@�Q��DID7������X����tJ��Ԁ9��5�f�*�۟3���� �0�wao�&!��j��>U<Eбڽq���9W�QhO�9d�I��\4�o�'j��~
�8/nf��TRo��2�T���)�ms#����^�&�u��3����o=yː+��$�h\h�{BF�7g�_�UT���?aɊ��Qܿ`���ٯ&Z�8�n\[g�d��Y��fFf�v�& <��%f�=o����ɩ�O�@w��!!���_���U� �2oI��y=nv���K��)_vd�/6�X��&��M4�q��o�CK	�YF 7�˭��$C�IE��h�0s���q�1�8=���Eߛ�p�R"ϛ�3�!�S��|W �1��Y8�rl�P#2�m+��x��ÞwRc˓3�n6��67)���h�#Sy��q`be]S�v����1;��^�^�0N^���(��}�7{s���^��Վ��jz�]�6m��:�5L%Z�6
��L��u�P\G	o���������s0��tg+�|Щ�ۺR`�I�MCC�=�P	�#�/�P
ܰ�a9=7�$�z�W,8 mLJ!�f6���M3ux<&����>���;�JOM%라ӝY����;�!�������|��4i�R(�
�B&�k�Ec}�8�c�`�z�;�>£$�(���3�h�x@yC?���u��/��B�r���Y�w*fp�	J	E�p0LAK�4E�u�?��jM;��d��ݪ�#K ��!j��D�jY����0�=�$�A3�um�f9}� .'L���O�+�5������b�_PR�TmR�Ѭ�V�O�V޸a����4�����t���<�,r�ʂ�{�$����]�d�+v�F������o����2z@��%h���쾐�D��X�>��z���a>�T����E���;B7�e��[	�������7yF��ƃ<:|y���3B�^�<�sC��������.�װ��Z�߲>
07{�U���H�ɉ���+��k+Rr�[��5A��s,��S��7��5I�lի�+Γ0�N�=�@Rc��HE�ɥo��!�5� �I�ڏ��G�H�����.��Ժ�;'!���G��ۏӯ,t�F��g�~��l�u�<$�V�)%��o���-z{�b|H���&� �4���l��f��R�"n�zxl�	�.���]"��� �<��`�	��F��蠃��l���'C�N���Й����e���ދ{_>�\j> x�<�DG�&w� G����f>��S������Z˻="jZ���� ��mJÅ��J�1�÷T�*�E&���,�5������k�A��{N�r�o�ˈ�4ʈ
�0M�xޤ$e(o��ڛڔqIr��y���
����|Aے�u=c[!��(���^�����G��U]E���t$�ҽQ6PiN�d�蜓��
�瘠�Z�o��!��[�	����g�FZ��_T{�1���|�
�qb��b�mk��,&d) ���:�A{A7Uy�&w��n�3D8��3FC6���n�
%g����b����PK1 �t"   #  PK  ў,J               126.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G.�EK��4�⡃yc�.�I��Þ���~n�I���'��_����G�d~�Kvc�߼������v�\9�,~Q�V'0��a+�o,-bLB3m���z���v�uA���l<�x��R]�N�?�5�kS���X�W�)f.�W���~�z���sկ��������p�����D����ɽ���[,�Tc��BU���E]80����Oy�.�תx:[֞�a�������r�[��]���Y��?�Þ��A}��o�t	ta��/�6��"9�B���W�3�pi_�����e�j��N�P|PTS�s����8���"b�P�/t߱x�ͅZ��K����^:���ǣ���7w����!:��^�����_�L=x;_�]�N��(�EMM�"���w���OlZ���r�p�B�o�7E��^v����9GK$�g׺_�7k�����"!�D]��܊]�����po5[�P�����{�Q/j�uί��}zWU���҄ʜ���²��y�X�t� ��;�FTM�]�5�Vh���]oJng�?��LtjJ����پ�u֡���6��N��4Y���0cQ>'�T�m�({��a��J���Qׯyl�|4�YY;a�+?m��9>�/�����Plw�3���	�n>�wj�ًl�r�kO;�U��U�k�\:t�(/�Ig��:.�Ω篃}����/*u+�<�}��2� ��ٍ�N��x]�:1�껋�[US%��t�[�*��mav�p��$#�u�w�t�i���t���e�R�?��3�	�h�~k���>0���k�Ƭ��ץ���\�p��+\&��	 PK�ݞ�    PK  ў,J               126.vec�e�Q�w������������
�؊�؊�`�`��νl���`�/�g"�,�(�d��yJS���K�(oWA�H%*S��T�:5R.j���kS��ԣ>hH����]�)�hNZҊִIE�6�h����Dg�Еn)�{��zOzћ>�����c`��A�`�0�ag#�
1�n�>�q�g��d��,��Mӧ3���b6s��<�1�n���E,f	KY�rV��Xi�J_�ֲ��l`#�l6�-le���Nv��=�e�9�Aq�}�G9�qNp�S���Yy��\�"��������unp�[��w����}���<�1Ox�3��YQ���y�[�;��|,����:�&�Gq��?������_�E�PK_�<j  �  PK  ў,J               127.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G.�EK��4�⡃yk�L+�oq84~|}�O6��v�B�o��-����+,�e����w�N�SN	tTt	`ă�]W�޲Ƞ�`�QCՃ����I���v��įᩍ5X�.�����Q|���L��/�BM�Lfu����g/[H�v����-����y�"%�/�j��H�{}㉿��MQ1��4V	��0���W^�O8�j����[�)��z�����u�c3����^s�G�jk�$���j�1��=%�ՐU$���ۙ�R�X�u��l.~�G7���xabl�~�'V��l��n�i��?7LOh�}���!��Y��`+�,�ҚKS2nN_\[�R:!���u��	�oZ�H�}W�c=�I�Z��,_�+��H >خ��vUn�;�v�ܻ�g���S|hE࿺���c�z>�a�	d�d� ig���C����\Xԥ�EȽ�{R�sCg���r�ݴS�9��S�n袝	��/�+�W�9A���ha�s�]/�m�{CHc���kd#M%'����m�ݺv��?��m��}>c��J���?�EW���8Gy���&���K�O�c����/~fҏ��N�`h�Ps�u���ܵ1-S�nG|�NJ�j�R)|X��v����N�/\o�35��̊���/�Vճs5�i*s=�g5����g�3�_de��%�,��)�z��H%�ʙS���6���2�}��U؂�L�7�o���{+r�$�;�j��k=��do�~�mӁS���a�㶣���WP���_�&��6���qܙ��7���xm�g��o�:B;��� PK{+8�    PK  ў,J               127.vec��Q�o������������
�؊�؊�`�`����a�7�=00'"�������)I)JS&壬]9�<�H%*S��TK)����kR��ԡ.��O��v���4�)�hNZ�*e�:�h�����@G:љ.)�k���ޝ����C_��B���1@� 3��c8#�Fڍ�G3���c<��$�7�n�>�iLg3��l�\̵���gY�b���e�8�ۭ�W��լa-�X���r���V����d���^����rqH�G9�qNp�SYQ��g8�9�s��\��xE^�׹�Mnq�;�߸+�q�<��ݼ'�)�x^��|�+^󆷼�}��G>���_��(�o����'��͟H� PK+Ҁ~h  �  PK  ў,J               128.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G.�EK��4�⡃y�F���6j�YZ`��_�Οzb>�S�����x��%�L���Y����Y^,4��Kc��Ƣ.|���E���e��­��6uS�m��z����ߑgf+'?���D\����
Gz�.e�|���laEj�Nj��J��5���#��?��-,|��]�`Şy��k��-:��R~�Ɔm�/u-d	t��eݶ��Z8��&1#�5�O�:�2&d���_���ޏ>��r���
��v�Kڱ��٬���b@c������� pL<����c�}�vO���J8����c�JO!�>�O�	WX�l�^�%�8����X4�k�.�X�7���3�2+�Y%+\�;������MS&x�n��(� j�"l����4�_-��1�ڢ.B�r���E}i)AZ;��ۙ_=�ß�K>��W�^(�ɵ�Oú�}]��6��D(���~���]k����J�+�f/�h�r��y�'V6N{}��o��C)O���渔[��P�wj���Fy��?��u�0����l犛�w\����e���%��r���_��W|�+�]\wU����V��%��"@O3����G�㲷;��#z������ks+�L��w��g-���4	���W������9*�9�jL�J�l��g���zOk��E_��Xe���>=`����g+/>s�%5+�U,��@W�QmkQ���;o��L�����䣩a�6�޺������2^�xY��8�7_f��PJ��)ɒ�4���?�=�1�a��J��<fx�p�hE򗥼m���*��I<��b��:������uZ�~����T��� PK猑��    PK  ў,J               128.vec��Q�o�^����[���ݭ�
�؊�؊�`�`�����a�7�f��LD���+G	J���)Cٔ�rv��
T���BU�Q=E԰��ע6u�K=�Ӏ�)E#��z�Ҍ洠%�h��h�E���ўt���BW�v���]�AOzћ>���S!��Q�`�0�ag��H�Q�h�0�q�g���&�Mѧ2���`&��͜���v���,`!�X���,���v+���b5kX�:ֳ�f���f���mlg;��n���}�� �\��9�Q�q����iy����<��%.��W�U�q��䖿궼��]y��<�!�x���煈�%�x�o�[��P��#����Fq|����!�����PK�`��g  �  PK  ў,J               129.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G.�EK��4�b�1���R�I�s��?;�������d��d��7�.z��u�ۻ*��Y7xU�/�j�S��)�����"��l���W[J�M�j�[�)������һ�y�+�Ŷ���"���f��#,4��k����b�.���ڌ�8%DO<��hw��5�%w�<gl���lg�j���>�Toi,�����+oMٗ����Ϸ��O�X����ݵyw����1��@��]���)�ڋ9}a�O���>�TZ�c(�n���W�U�强�W��a�ܰhgg��E�&i:��e��*�L���Uo���[�K?�I9x�����Sj��K�-�}lr��g�J�����*�t�M=z�V�K���i/u%��2�å��|ض撻�	��3�v���l~�z��l��ڠ�^�EM!��{���z�|&��;ѽ�H�O"��cw~$��{�sUk��&G�s;g��N������ַW�
I"�C۬c���ݨ`x�S���y�$�aQ��\�p�̛C)�tc�\���d������z�`�a�����_v=�~/�6��ԏ�N]+54u1�÷>枺�=��Ӏ�>���@�%�u]��&���°���[�=5*Z���ڑ��[.�=�M�̽�԰�e��slI��O��}��f`T�nrn�?�}�D>��y�n����f�J��]�y��Pf���I]Ex�m�#��k���,�~"�F����y3r?ʾz,����0��;)�j];g.[i���w*eDۺ?�K4���R|2�s�'�7�6�֒=#�d`|��AՉ���>��[]��%@p"���ٻ�Qj��]t����?��(�ߣ�{�С�/��r�ν����ξ���{��9f��@/��K{as&���%�u���K)~��u���M PK��A�;  N  PK  ў,J               129.vec�U�Ua�ѹ�n����[�݊���`��؊��
�`+�j������VD���/G	J���)Cٔ�r��v*R��T�*ը�R��մkQ�:ԥ�i@C]#]c�	MiFsZВV�NY��"���hO:҉�t�k��壻݃���7}�K?��B��Q�`�0�ag�n�n�=�1�e��D&i&�S��4�3���bv���\{�Y�B��%,MűL��^�JV��5�e���F6��-le���Nv��=�e��\pr���(�8�	os�=�i�p�s��5���\�*׸�nr++����r��<�!�x����3�9/x�+^󆷅B�s��|��K�����������w�PK|n `  �  PK  ў,J               130.i��eX���nWRz��%�SXBZ��E��niXB@�A���i����%���?��s��}q��r�9�|Ιs�;���ϕ��h�  ��<.d���8�X�888xx���dD��T$�@2:j=5--37+'���M����W@@ �**!����_��?�����RQ�1�2��?�c�M
����@'F� F{�����B�o�CC��������'x
h|@G��@������|��?���X$���ؤ�f8L.d|A�\\�Lm7���	3��`<|��T�,/Y��!�B�"�b�o�����u`�z����V�ml��?yxzy��|����5)�[JjZ^~AaQqIiY]}CcSsKk�Ϟ޾������ٹ��ť�ͭ�?;�ݽ�ӳ��W�7���B`��O�?r?q�cbb`�����?ĘX���$Қ8f.�L|A�d2���n<0��	��I|
f������7��X������\K B���� @'~;y+6�4��T��,B8C�:{���*�Zu� Y��:�XtJ}JE��3�!A�tʄ[��Oj[dUYfiH�l;=�h�R��z�ͪA�HB�c5�ʲ�_Zv�ެA���š�@�@S8��t�-f���"6���ɧ�HR�x�{��Z{d����n����uԤ{;1���}q}�}�ԡ�[٩�����y������Vb����Mc���t�tX�����u�P[aX79���c���L��ʽ�rf��f5�iI岝���"H�kqh�#\���r��g�V��������qWA*N6�z���^Zu�[I>�s��Z�j�3&kH��nA_�&�%&GO�jtv�7�33�g5�GV����=p��y��=�0Bg�li�%a�-A�tI�CO9�V �o	�Z)n��� ��]ĺ��:}�_���yj}}@t�$g����q#��(�s~���lt�]��zGE���^�gi?�jt;YSr��.ee�M��qr�6ضb�N����i��ǣHՌ�+O�m��ϩz<�1�l��4v&��n9q��l,�	��|�%�`�(�#�\"�ޔ���?�uT߷.Sdb�ӤF�����@>;x���pm&�6Չ�c�-������S�`�B����ۯhh�Ev/�?�k����p蓑g�3�0wJnj8�o�hKF�A�����6\�B�?2�?{Q�ZA�s���oO�����:�j-���XȞks�9/5~�Za��8�)O\�ۺT�`��n�4�9g�l�SrAG��m�BnQ�q�+�y�H�12d�eG�:嫫�/Wn��^�5P�с�a�o�&m�4�/=U#ŶJ����x:㜣���>�IӍ�4Ќ��2�DՌH��G�a�|������]Шn�Ԍ�����췧rw�
�|�?��Z[i�}}�	#�Ƭv��U�cx��ֺ���ҿ2Y��	�������n�� &�R���Z��b��~�\���O��M�G-I�ؚ���r�(o#~�MB���B���u�_���W��烾�d\�XZ\�#�۶"�?ZM�|������O�����if �pI>y[�2+����4����T���Ye'��ف��}�����YE�m�����^�*6�woL�Uy��1�]�)_��t�������F$�sUԽ�����W�����XZ)t��j��$l]�J�_�vyXZI��݌��ޞ@��f��oo���M.{Gj��۪fM�?nv�|KF|R���� �Bn��-Z�$�*"SG>��-fM��Akg���;�N�Bm��s����W)S��ȿ+
S?��B��bx���)���Tm��a��6����'����G�Ŧz��bXeMʟ4<LK/=js@< ��D�S10^�>偃��~�u��r����[wTg%ỷ���آ8��X�S��5٢W�V�e�;��>�Fb1�z�$ ��슍�_���=�;�=Ev٫7}�v�n��ۖ �?AO��WP��
oأ�ځx�.0���ȁ*sĺ��^s��(���2TjUm���h����Z��ܜ�Jj�~9X%4�Y�\ K� ��v��聢v�������%��� Dj
�WE��˩�9W�;�)Ac\���5���&&>�՞�7�~!*ԣ��끭S[����*>�vk+��,�Һ�-tB-q����Y���S:���Z��I�]�!�F��1	SʃCv�p5�u����m���7�y�#V��������w�G��߽�X]��,�)Hi��e�/j���_�QN�J8Uq�H��f��V�5�.k�&�uB�8J�����*_��݊�;q��ok���W�J(������"�g�N-���0�+Iu��@wZ��o�8�@!8��#Vc��tޠU��n�(�U*�?����XV� ;0�z���q}ɉj`U,} M_���0k���3tK���`�����V-w�p���..Ӽ8�p�AkI<V�k�\��ݤ���T�؛�3"��c��k��R3�D��Э����G���/-�!p�-�����T�K{V���fK���!;�G ��-��#@��(\"z��ͪjQ��s9(#�}x��g�R���w���W����+���<���~�7��e�Őj}R��ע���.���	��m����@�a��zV�=r��}�q��?]�3��U~TlRy$�MS�<gT�L8��[$��
Sےa�u��>n�`
��+ʦ)�������b��4{Dkے��_�����i��4�v�׫fj��f�5j�r=/��+^y���d��%��d�� cn�r�Л,������}Nm��� ��֬�N]�OP��}�S#f�>�%r��!�ٯFv��!,5k��	ү��"�31�� �j�vLcA����*��h~G��@�G@,*�}\�]3v�8y�2�j22qܧR�(����;3b��~��]'��7[н�����o�BN?�Ip�=Z0�/����%m��������b�BT������w�Q��G@A��d�-B��R�ܫJ{~#���v��C�h�sh�����B��g��'�i�S�І�z~l;p�?(�ϊ��HJZ�u������Z���Յ����R�2o��G�0B�02�Ai��b�2K�Ƅt�ҷ��?:Ք�C sk���#
-y]2�@�T(x��[/E�5=b�go�1�����-�/w��u }��T#a��~�p�iӰ]�t���Q#���q�odW	���o*�w��A�;�����{_P��؊��Y0���"j�I�������i��ɍ�p������F�9]���u,}�Z�F������(����1����w �i��j��#�KO��"�ƒ9�E��)�{�Y�T����&�g��S+R���_�-��xdl,,S��px��j��@d�iΔf��"У6�B׹0o�,�&�t�E������&�G��@�#���}*����!0-<V���#`1��m?�#��|l9\�����S��z�#��~��(���:���i]ng�R�Z>�ͦ�u���AB�x$��˵D�
~�u%�'��ND�[�7$�]����Q���+6��M���#��>�����V�Ѣ=d��7ӥ��� �a��Ѻ�KH��_�|JUܲ�TMBP��N>q���Ϩ�ן�z~�}	���O_m�v�/6��ژ��{9{���ÅMK���j��e>����i��\yǦF_�V���{]Nɂ�����"��K���y���s2y�7�R(I1
Cm>E��q#������߅�^#4>>�z�pR�nv�(9�v�N4Vݸ��.o&�F��W�p,�7�p^婾C�����#����2���w(���71���.:^wSF_��I!"ʔ������r��k��UXٙ������S�o�W��-p����������)���PR�C"�tC'�ꈞR�3F��'Ly�T2�~�+�n��'W��/�����q�82C<T��wx��Hnm�S��ddt�[N;њcB��2����lH��K6�C�#�}Lэ�i�}���;i��h�%3P�� `F���m$}Sj�P�B�����n�$i�_d�S�����-��/*n������=�*u�Ư��Ns�^��b�/T�7A�ԗ)Q���ac}ǭv�怒'����C��-��C.dr_c���ݘ����zb4
��'�^�SQ=(��˄�k��\�Z�邈b��G��[0�p����v�������kD�ry�i�/��#��Xu́={�H<�#�ޣ�+`���W��m0�f��6n�<߃��剸E�r,��������w���eq��
7QA��gFi�B;��	5���V�WKd��5�h'S=p�{
ck1��l��c����G[�(`�厬g/��T"ݾ��f�O�-��'�X.Թ�)��rSפ���kH��T��V�Q��c�L�R�\[1"��b2y3|Kf1�)���xywiAs�f^t�v^v���E�e�ɼе�G��XvRW.�
`�J���X��;��2��ɨ����g{|�-a���ӽ�y�Yi�U��4�A>|���at��Rj�ti	��nI�b~$z����$���ytAghM�E�i�E.b�����I�|�Q��s��N%�~*�*�l�u3�ɜ�^^_"~>�����iJ����_�x����q�7��4��# ����Ɍy{J�x����o��Ӕ���3[A�
�L;��z��-Ҩ9y�];���n�DɖAX���#CC���O�G�5�o��!ŧ��ζ�&2�h���[�%���/�v� �������w\��t�TkR��P�g��Xn�]��+��3Wc�T��1��Qq��͠�G�z,�Z\�u<����.���z;V�A�PT����k��MK�1�7&����F������s������r��������{�oT�I}{� +~�3C~O�5��d��,Iw�
��`���U��Y˙@X1�$�:cj���{�R�$�p4=A����`��hD�ߡ+T�2ؽեK��8�m����dQ� �*ٯ�>:Q����/zt��c6����v�Ƚ�c��;�s�8k��^ W��t}Ԉ7��8�r� �EP.9�ѹ�����{�G@P��Lj 9���~�h�nǣJ��p��~B��BZj�ˢ��Y�O��A�r�Z�z���ǒm÷~OYX"��=DI���?��i���ڼ&�hL���0K���M}y�&�D"T�(H�5 ��+�n=�$V�*4�ܒ�l��Pr8a�VuÖ��%H]
��W�<�4�x"�N�cU-IR��;-��3���`�)�{�!D
�L���������`Ajѿ>!�	U�%mF6m���m9����"��T�Ծ;2��_V���j��uQ����R}�v���a�׾���j��]��7� d5�#�Pq�?�ߗ}�:TF����5~��5QR�p�_����[��w2S�M�� ��>tQ��)��zVԁ>�~(I��JD/�1pqI^�y벊C�Ġ�]�PU�F+����MWw?��8���JN:/�u�5z��?�0\�< ����_�v�Ml���� �����𷳘��H&������aL� wA�4ntt{\˅#����{��^HH�Uv��2�k�W�w�G�sNoP2?�7��ku.���F��Q̈́�hL42Fc��Ǯ���Mڕ�Jր��e�B��/E�yČV�=3�<�P��7$:Q1�a[+�61�J�V������ �ӛ�����X�y�юL��),�r�<�y4�x�i�kEXYA��uC4��̾���[�o�}NSJ�l����{�ʋ�-�l�y�WbY�	F �Ұ�]��sW'�1��!�`��'�φ�eр*JZL��7��{}��ʰl�0S���ĸ�>W�������9�1���At�^ �Ea�s����4ن;��{L��>c�ԝ���}E�'��v����'O���l6�5�H��O��"}6��ҁ�FXx��V{���p���k�|e4#N;���U_�ª���?/&�;:�/F�@���]Q�+�y�#ks��F��oo�?���}�qK�����>G��w?G�jKnG?�f�]�'��MH�\�8^�O_��i�պ*��o�fMF�e	��k�ZIi\�G˘*Y���Ӄ�i�1\�"���Dtr:��>�p�>���>G[���~�H+Ht�Xӆqr�ӂ�5ֵ�\�9�32�'�w��~�K�[�K��\&�8���̿!��?���ٗU��{�����;��!��/���w��.�3�7s.�d�B�,��Q9[%���ȵ�a�O�Wa�J��	N��g�l=Fm���D�Ii,ܗ�����@򯃡�]!�k�8피�L˘R���.�|묜o�3tz�2��	�ɚ�ε��u���!+T�Ӝ�hi�L<C��pֶ��+�t�~֢� �PUbwh�V�f�y��I�员��.����%�Q�4��:튙�mȳg����q3��7�tݴ%�=A�F��Ĉ�Ŕ����������2}�	a�u�9R8{�M".���T\�Ϊ�ȹJo��"�݅^9O�5�e�af���zt�P@[C�L���}�P�W�e�ɖ������H�NPV�������͡�-�g�����V�Ҫ�>;��B����-��$�VM�%�8���?$�d���[@d��M����{��'c����� �{'�Iiܸ)��X�`��&��k&x*2��Q�1`��
�����@��zNW���v���y�2R���d�� Bh���T켁���𗉬s�$B�T�M��;)�3�>W��⯊����8�/��8��.D��%_����NQ���QmE���t����ao���.F�7�~��	t���
p�,jc_hJ}{�+z4Ƒ�B�u�Y �f���I���hX����5H��S-X�.�Ml X�Kԟ�Y��������e�d���w�vP.!?���������P��E̾o�,eZv�:��J��=	�b��ֆT��c>~Kސd�s����?	T�-8v>�3ktуW%�?�<S��}R�ʢW&R��/���s;@a=9U�m�$��	goP�V%��hdc1_�كE�<��X��eo�Km�&�;C(���z�|5p^4�Hǆ"�����r��>)s�0�ǫS�E��Wo����~�X��-ӔQ]�#>x#nF�v�Lܯꑢp�8D�xW^N��0�q�(e^��0��}YfP=�$�GY�z��R�ۆ��W���x�m�A�:�>&��q�j,��#����8���Jz���pD%sM���]��+������F���P��F�v��o�i�ʋ�QBc� � @�%Q��oY��Q >eg��hB:����~N���Yp����|���/e����u~S����� �${ŦbΦ>��z�i6�1���Jt�k�Mx���W�ǁA��8ta����E2���H|�م��{��q[���� ҅~��1��TNҕ��Ж����E�����
��Ʊ���E��'9mA�Cw��NOt�`�J���\�I��n����`M*fM5n��ou)z�!|=/�-�-�N5õ3�5��l��k7㎝7����a��k?�i5z�ض%ƩA�2�Ep�"�c{�i�.�V�<����^{1��ʋ���
�A���h]��?�ȄBx�1�V���w&)/������3�V"S����" ih?�v>�q����IP�A���"3�s��s/���|�{q�\� #������/-〃�Bw��̛=��As�e���EB+��DiQo�f��h���ټ�ME����0���b�S�us���n��{I�w�����B��M9226����{���.E�Sd�h1w�����٨0,F�Ym����4to��&g��<Y-�ܒ����k��e�X��t��L�)����`?ܯ�n](آ�P�'uA���1�aʵ.�U=o��G����q�Rlb�~�(�x�笷�!���u���m��#@y>���۪e��~]y4#G�V����+�)��#������=}�6|��'��8�qM̘��v��Ә~n�g�1$�*�ε����>x9��U���
�7%<13M�R[D�bP�
Y]��8��]/��2��~B��ni7��+q]�t��$�"t	V��{߫���{Ȳ{+�f���G�
���6�"Ӕ��+U4�fh�3����}��F;�L����Jz`�g7������'q��ն1?R"ʜ����pЛc��igx��g,�P�b�A	W�Ҹs�!�ME
���'�s�QO����A�m�pf����;��d�Î\at5x����$�!TR�78�7y�����\X��%m:����&��sջ9y��������Yf�fW���V�S�,�)j��p����d�(�|��.�KՓ����!���A6C-+Mz��FW�2��ʻ�S�d����DלIPTf����o.�5H��L	^d�΂W�yZ�3i�$�#�S9�c�llly��d3�6
�2�v�D��n�Զe�����F;h��a;�׎�<�fmW"����'���/A3:��vM��ܥʶ�:S@��+�S'�aS�|x��<ؾ�׺�$=`�6$Nl��䆿M�i�7���m��Lб�{a'��fZmv6�Z����w����h��맠L���]�mm�l�O]��oG�Q�̢[.%r�H>ᙴh�����PKh�X"  �"  PK  ў,J               131.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G.�EK��4�b�1�����"����)�ϔ��4����O?㩶����tƲ����p��w�kS���;sui,�ta�#fܺR4Y���w׻o�z�QO��$�z���_�3(����㕞�H:0{e�K�%�7����~�ܻ�}��8-n���J�-�(��`�;<������g����*����M$Е.��}���]n�C'�i<��+\�?C���'��pRj��Q��G;,�~�W�H�_}F-�����mO��iw޷��p���	��mP��r�����+�����X�t.�j�n��+-^|�U=����Q*��-���X�������'�y�S���}�Y�7�EwE}%�ٱ��n�̍{�=�������nz�ǼG�����W'N��|�գ�-���nX�U}Q�f>���˚�Dѵ�W�;�q�-~�2������wZ��|��|ҝ�ߖ�Yŭ�x���%w�]��\�H1?�H�ǆE]x0s�!7�3�����'�L�}�u��e7_�Lޜ���.D�����k�nL�mtѤ&A��/x����齋DD�s�//��&���wk�`]�|&��Osmg���e77�H��Z�ubq�$�Ӫ'�a�+�T�._3���o�.�0����j�޽�&9��_�}�=����5gO��6����������X.��}�������w?��:�����|��)	��8,O�����Ug�+��[���E��W�{�aa;���q)N=��lqv�+�x��z��u��u�&�{��Q�P��z�Ɩ���k�z��s��1A�sf���q�>�k�SY�}!�Ve��y¹�d����9��X���WZg�mZ�+�(�;�w�s��$��7PK��#�*  >  PK  ў,J               131.vec�e��A��=�cwwwww7vw؂-�b+�b+؂����s/�a�7��6�e���(EyJS���K�(oWA�H%*S��T�:5R��v���ԡ.��O�(Ec�&zS�ќ���i�"�f���t�#��L��ͮ{��zOzћ>����
1�n�>�!e��HFٍ���e��D&1�)6S�4�3���b6s����g7__�B��%,e�Sq��[��b5kX�:ֳ��lb3[��6�����b7{��>�s��Y.���(�8�	Nr�ۜ�g8�9�s��\��y�k\�7��m�d%qW��>x�#�<�y�8^ȗ���F����� ?���ȯ)ߢ$�G�6?�/~󇿑�PK��F�c  �  PK  ў,J               132.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G.�EK��4�b�1�Δ�y��+M�vu�}m%�����ʞ�Y_��l6oѹK�ߴ��K���x��;��W�Ԯ�lo�/��FNtv,�^��Λz�y��`����*<q��9!SEU��+��B���K͘r��Q�E�������q���Ta�qi�;P����`SV���-�q�3Z��׼���?�t.9W<窚��.�E��"��8���z�	�.��i�W�d�nzd�����Vo�e�y���?�Jf�����cL������y�պQ���Q�؞�V�_�wk^_W�_�sG�Җ_~m�)�oN�c�;�L���H`�G���x���Y\\�l�0~�z�zp�����$��Q�����r]����&�7�wlw	fXԥ�3/�~�S���Ͷ	酎���_��Ur������1/o����BOi�u�ލ�Us����4�8D �������MWH^��	��O�]g��m���%V�o���/|λzzޒ�bq��Tى"�.
lߘץ�$O��a��أƖ=�54�1�ў���n뵊c�!�j�B9��2������U�����ԺRCcQ>|�r���U��1r_~�S7coO�Cߒ{F��v3/�!?imѓ9��e��g�k��Ǵ��?���fF7�M=������{���g�������>�OlO[v���jv�<l�׿�7ݩ������Ư�廥�lv	��O���ۮ>o�L����?:Na�uoݷ�������[1��oziq�R�c7X���P���3�3k\/.9��(�w�*IƉ�v�>s�q� �X`�K
�˯��\j蓙:�_����G����y���35&�]�!���;�%ֱ����������@WE|H4�zY��䀮j��u&�T��� PKǅ�u  3  PK  ў,J               132.vec�e�Q�w�������z�V��.�[l�Vl�V�[��S�����a-؋=f"�,�?9�(E�Ҕ�,�R>��U�+R��T�*ըN����]-�6u�K=�Ӏ�4r_c�&zS�ќ���i�"�f���t�#��L��ͮ{V=����7}�K?�3 b`��A�`��P�1��LY����a,��&2��6S�T�1��d��㮹v���,`!�X���,���v+���b5kX�:ֳ��lb3[��6�����b7{��>�s�;�C�G9�qNpҷ9%Os����<�ȥ,���r����&�����y�{��y�{,��g�B<�/x�+������{���|�3_R.�FI|��m~ȟ��7"�PK��bUf  �  PK  ў,J               133.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=�G.�EK��4�b�1���-�Ek���]���}�F�����i��6�����䊾�-:�n�7��+b���_+Lfɵ�R�@GW� F:b�g�km�zv������SW�k�?���:)A���F�Ԏ����M�J/�����m/gv:TW���n���.qL����]��\�s���[�7e�>�nѶi�����V�-��4p`���nMO�o�u\�g����1����-�u���U�.A�jN�<�Ӓ���-4���ץ��ֵnON?�sRJ��S��$M�lm���͝s�<���A��Ԇ+��w�y�{�´.��*��p��[OwW��^<�j_�dU��<F��ȴ\���Wg�y-��ϠՓ<9�Y������5K��]`�J|���m����[�I�\�9f�?����x�d��%��:o�9�j�Y)�����m"qK����:�����=�b�%�V�$+<���X��FR|��_o���}�{�չ�o��ɽ���W�sٴ�ֽ�S]�p3omՇ�ګ��T�P���a]⾏���?����<�o�;�'����ݘ�ۊ��d�c�3���c3p8(�Zf�����[��-����_��j��gz���nru�=5Y�Kc�t9�3q��Ќ�)�N7�_�R7�����F�+���.x��� �����6�p�`��X}��F�;_bM��	F_��9-�p�		��\�2��?e���ﺙ�=.����J�U�=�H�����>ד����0�a����4���I�L�;=LO�X|"�hA�i���ޕ��b��
y���0�hJ�P��I&��vܐ�����mύ�ʵ�eӟݓ�x"ݩw`KBzף�l�/�j��,��X�/����ꏜ3Kz*���">��?�#�a����G}�N�>��ۻ_�Zf[����߇ث
n��v	�ta����g��gؒ�诮w�� �S��M PK�Ê�e  p  PK  ў,J               133.vec�e�a�=��cwwww�[����l�[�l�l��O����a-؋�2�e��)"G1yJQ�2�M�(gW^�@E*Q�*T��S�v5�ZԦu�G}����5֛Дf4�-iE��&+��z;�Ӂ�t�3]�j�-�Ew�=�Eo�З~�O���c�>�3��c8#R#�F��X�1�	Ld��d9��Lc:3��,f��1�n�>��,`!�X���߱�n�����b5kX�:ֳ��lb3[��6�����b7{��>�g�q@��9�Q�q���Iy�Ӝ�,�8�.�\����U�q��������]�q���#�P����y��R��5o���w����r�9�ėH�����~�+�?PK�pe�c  �  PK  ў,J               134.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=Ç_��0ui,Ťc� ���w�ui��IO�9(�����/�M8Y���b�9���ͅk�߽�S����뭯����j���oRXԥ١���������Mb�κ#���Ң��.�l�'�,!��c��<��1��_ͼ_�I�t���})z�|~o��?�C�M��:O��=NǪכΜqZħ�^�����w��'0���zgJ�H�+>\u��9���5\-�_�Bu�:%?����nGM{����aH����sF����5����˚���u�-'ω���`���3s��v�/k�;w}��'[)�v����EN���/����Nri,j��������jo�ӵ��g���c;V��ޫh�۞t�?C���E�e9��&�P�(�bQWA��)_^��ʓ>�UTx��ސ_�����^���G��vW|O��������Wzz���yo2u[�Ӽ]E�%]E�`ƫ?V����U�։Q��o/t=~�wcQ|��X���^�2�E�VY6��ROUk��/`��lZG�β.�%���HRo�u�O�`�+��~���{���+�ZV�����{���9Nw��.�^haq�?�����ŭ#��_��-]��������b��a-�5�`�A�w�o��o���|����' l��?c[ԑ	nG	X�>��7{��'�n�Ѯ>r}���r�����-���2��k��r[m���ڏ&������F��>��Q-M�^塷�-�/W۫����G�C������^W�8�?Coe˻�]SO<�	Z��}g0K/Xԥ��3=�L��{K��[QBv5�����;��=�ZvRe����J�Vu�/�>��7/t��Y����ϛ�ϟ72�p=���2W���g*���ڿ�\���]�mS�>宒K�s�h�{�e���uK������Ҹ�?���;�3]�6��v�y�8���rޖ�S][EXq`�ˉ�w�
,��l�֑��7PK��K�m    PK  ў,J               134.vec҅�Q���|vw���k���`��؊�`�`+���C����.�a"�,�?��Q�<�H%*�|T���W�:5�I-jS��)E=��z҈�4�)�h�v-�V���6����":f��w�]�FwzГ^v���G�K?�3��b0CR!�:o�>�bF0�Q�fcS%v�z��&2��L��*�1��d�����7������E,f	KY�rw[a�R_�jְ�u�g��f���mlg;��n���}�� �\��9�Q�q���oyZ��,�8�.r��6W�U�q��䖿鶼�]�q�<��y�S�
�\��%�x���������g��\|���n�C�����PK�FO^  �  PK  ў,J               135.i��g8@��U��YV�(A��Y%z�$D'D�Յ`�N��{O� V_a� z���z=�uʗ��s�ǹ���73w������\UQE�� `=��@��>>>�#Bbjb""b:J*2jz0#=��������q�pr��		��ŤD$y���11-		��3�3��g��P<����X@
��^ �a��X�m��aX�@\<�G�DM� l, �����0�0����|�/�G�c���F-��{�"W��F��!��;���Oh��ٞ�spr	A�ED���_)(*)�����6������wp���������9*:!1)9%5-=#���������������������W�`p|=95=3�gyeum}csk{�����������?\X  ����#�6�?\X�>�q���}ƏG)��o�F�,��Z�W���EP����o�ǬB�lG�A�o��;���/������ ��X�� @���K詩>�o!̚��5��(�A���d��m�LTQ
G�G"*���O���3]�-7̟�ӤQ���#JKc�<�@�B��-i��@?�^�f{6p�U {4/��gǤ��f����Ԧ� V@[*\��{�*1�"�z��QC;V��4����d�H�RH�i��B�GUP��く��u���z��Su�v�͂^������g��I��綕wH�����/>%�*&:M!������v�_9����u�~�d�f��|�����ɷy��hi��WQ�Y=�?�6��~�o��g?��x�ͭ�t�a�Ԗ��>ʍ7�18h�Ѥ��m#I	�M�ؑР��s�_���{��ԧ͞��q�<̚⬊������@Nk����¹@u/�}�\"�pV6E���n!&���uZEG�5�'��!���5ب ���)8��捨���bw�B�{ m������/{k�'�2_c�_��g�S��)ߖ�n��"gv�e��s��?�r��~iL�.�-���фrmV8�{�����:O 
����8����A��sz��hf�rGi�@�Ft��6#��\h�|��#��Q�Ӈ�__��o?I�$V8�$!\%�ia&y�� ��=�#�����v���-�J^~��͛��:�����o� [���ݣ%zs�*�����m��t�e�N�~�!���a
$���\��J��c��y�U]b��j;�,D0�Swh�jRt�`!�Zv>3���K���*s$�r;.���R PB���{V�f��Ny�����4	nB3���{@���xI)�<9
7�+%|��;+�i�y{p��*[��4���apH	Zu��^�yF��ڬ�yB(U��Xg��K6^���|�#K���M^����$����Ћp�ϻ��g�Ȟ�k:IYa!����T�3�f���:<��h07{Ez�P��!]��0N7�Y�������TNV�w!/��� ݿf��t�M״�5��t�+��}0'^������=	�m�����'j��~9U�����(�}<��]���-���f�56�Zn)�Ζ��f��������o:�E(���f�j���P�,�m� I+V9D��~��0+���m!�)�����j�U��kb�<���-)��/1wS�o�:�.�=��&�j���V
9��\ܑ�j�%$���+��Ρg���YE=�xЬ� d?�AT�m�+[V�&�/]"l��UhN��!�L�/|�픰`kr��wR��Y�_�5A2�,�K<�Ұ�{��o�E��|����̶����}v���2W� om�~�yD��4Ϝ�;��a�a.lݰ�Ӟ���ú���Hbkֽ�/�16��z�GN
�**I/�i�3���dl\}	�r�eN�r��|,�BL�9���V�7z���3�]�>K=B��R��Ye���~VV����6�L!�h0%��a��`��!n��l4��,�rS�l�#y8Vuן��8	G| �����:�ٱx��d�䲦�f&꫎}+�8�'rNC����M}�@�n��z�O�U� r���,�i�����92LΑ�E�PZ����w����������j�ޭ��A�Go�6��3�x��8���K��;�$�@jl��F:�m��8�>��~�_`��T��}�B��:�����L�(�r
�F�.�0y������+�ʊ��B'���)7��R��S��#��V4��GJA�?i=K�6�׮TN�t}�Sx����E��zn��tPS�d���e^�rx�"C��me��R(�y����p>zV@��:?!��^�msJ`t䦺ț%���̒P��6$�T�k+��³����o�J�de��Q�K:�T	���IMU_�����韉���
-Y�gdp�'�`D��#��2^���~����j��������C���m�V��xv4.�|�9<TX��8꣢��&������h��1�5+���gx�Qc�Ǟ�׋�Η�.�|A��K�t��fa-r<�+�Uܫ��d� �(���D�@�-W���`�i��n���r�3�1y��&WjW��D�������c+�8�`�'=
���5���,��!��z��CM�����-����pgv��k\��ʙ���;��]�SÀ|�,��ͻ�z�k���.�t���}"a4GU��}��V����]�=�M�i�ߏ�G�w��3�C�w������x%����aXwI�� ������+<5>|?�Xr���:d�Sq��R!|��o���C*�:��*\a�l&ޝ���1mR��� �C`�q�I����ŧ��[E�؀��$���usp��+Yј�}O��Q�j���O�g=VC��R����:�nL��m?p�GC�w��/o;G�阷�uP��������>����<��0{�@�����P3N7�j[���1��M��-�X�=����G�hyF�t?��_�jB�>4�4C�=Y����-hI�=����y�6�&���	0���������Ō�iZ�ɷm�&]�2����e$s�T���:w��*V�N��)t<� 0��	F�_OT�ߪT��wW�
4������9]<�0�Xg7�FW�qp�����\��O��8�TO��Պ;S{�r������)\p����uR�%���V�ԃN��*>��D�s��
;���4����rx ��L������J�{�婏��ET�a��p	N��EE��$��$`�O�i�vS�z���Ԗ�ߔ|hí�D���DO)�O���4����IR�,Wp������,�nd�`P|�<sȽ֬��Q�wLʏ���
�B�#i%���2a&�+�p�L�Q*�1`4}�s�����J�Gђg=��D�ab�{����
d��0ў� �P;,v�!l�?����w,d��jK��n�BM�L�DĨ?�k���#�!^Ho�\��z�̛��uR�ck|;5�"\C���F@l���˩c�~���!0KsJҽM|�� %��� P襳坂�����[ �tR���;���~�b��6��iA�D���<�j���J_��>����5��i򸂼�\��.��h{DH�梊6ߪ��ϡ.qy���2Ukܪu�j� 2���JNDsq��
�C�����tқ9����O����+��^�A�M~����׼�x @�@��>�}��u��5c�����U.��\��u�Jr
�[�q��s
�g`a�	�Ɉ��?�Yf�eAԨT}�	��m��z��P�,�`�R�T}���Տ'MO(v<�?�W�����7�@{�G�]g�� ���~�k����L����{�l�� �g�zml_$�=�B�@C2���q�,���=ܝ_���?#�W��;��w�'�'H����.Z鬒�i}����X-r9g۔s#��+��?��-S�}A�#P5��'� >5,n�i{��7gj3׮�IJd�>�&��PJ�Р���ʊ�R=rV�vGt�@m5���w�:��;GĶ�Iº�fp2XF�ֻ���}D�p���E�f�`S�5l<	�Q c�5�pX(0˅��=c�ߨ�1u�������I�0XzT��ڎ|Zp�5RN��-7����WnS�&����o����pJ�Q/��'���)0�iQi��������;~!^��m�D`�Do��I�o	ͫ~�1�aY�,��+.�~�_�3�L��,���W�*uB�E��)Č�V�}۲B����ޞ�Y6�_��em��k�<�{4	������� k�o+D4ۥm+�����?W	��[/�~�>�T��6X����FL(wd��P���"H=K[�� sKğ����0�A�K���]����.bu����[X����c�މ��JW@��3^��#��2�H�Yre���'w��7��E!&�q��<�z~�UP;�:�N��;����Ȝ���4� ��fX"��{v'�����i6�a�N��:xu�\�C'oȑ���uM([Ć�zs�˓�ʐAZ�6~4,o.]Z�򧴴���и����ǚ�2Z�C't�X+��3�e<J�yQ!ДM1X����Z���<BwN/�4]ʉup��j�������l�7>�=�<���*���h�>�LU\'��$	R?�~�m�auq��t�b)ɽ���e��i��lq���� �-�Ѯ���}������/���5��z�\"�i���Ed���S��q���*�'��BS��P�Y/2�� ��M�}=�����!G�+2����в���(��'j1��0�d%g����Գ��X�sw%��Ҡ̰=�����}�"�c�5U�s��w���c���Z���ZAt/� 

!9��yi$��F�%,Վ��:3����d��P�y����L4�qU��0>'��iz�c[�zW�[�G�	��o}xR|J;}U�x���[CG���R柌=�WS���暕|�)�S�����l����]�rr���k�w��G�3�����%�N���-&�NjC� �_�Vm81d./,C�r
�35`d�fL��,0�q��py�v�§��~V�M8�@r���<���<�z�v���,��B�����;@��5���I��J���/>�|ήż��7A$��Oo�S����(P�b�����Z$%�Y}K���h0:�U�7�A�������Ƶ���C?�~+������ɵ��B�U�?��-�j_������y����U��ɞ����*�7�gmX�Un�ӫ��)~�9���%����
x�[�L�Ȫà�c�R�X��?��n��X	5w��"uyd��'i��?Sh#����)�z�+��ht-�EJi�o1��v��f�ax(���A�O5Y^�֫�Ly��ھ��.�҈-��E�$O
�l�-��J�:dq�L�us�uW��˹ʿ���@�?�v��9��/:\��\��zu8r�Z)4�S�Y���i:�]���6����0��uƔk	����c�iv;+*�3�ג�g"B���/B�P8q��dբ�m}�B�c�>Y�k`hFFo:�تN�
�1<�e- ���m��z��Z������K�l�ꥊ�MlZ��q��ǅk`ǐts�0�մ2���oj�e�co���
�(������/L��MI�����K�"��
;�l[���-5���O1/C�b��������츒m��s Y��]HD^N�5��5���q��wW�v�A>�x�V9ۆa#jQ�B[�WI*�6qPu}o0k�,��j��I��/���ϣ#���w���T!A��<�ܴMM���_�"�+�j� �m[��˘[���k�&���^�n�S�PӿC�C�r;�D�;��CT�'. ��F�A���i�W~�	�+��lw�m7O��5Y?Ty_��8�aεm��'�a�]c�~����c_y� m?^u���������07V?�E�������Yn�zMQ��iv���(�\��e��!�NG.8��+�:.H9�M��&��y����3������(�ڍ�)A�"��V҉|u�,��H��bu̑�ІW�l��RQ��w�����1� *�M&;P1��^�^� )z���eL%(�1�\�+���kT�\�,�!4a\�r�{(�.����`+�6h��\����w��9�|S���7�1���7�J�?�Ak}�v���44�mQ �T�X[�z�����5�5&Ԯz�(���sy�,17L����Ӣܱ	�\�o������?�BK����P�E�P|�춼W)�-��*���*��;����4mmu�n�*}f���6\=a�v@ux��/4f��ɗ-Dlg&F����E�D�{�S4�'�4m�n�~!���N�7���j�~�к�s],�6��L�]c�E�0a��p��,��Y*!�� ��{�|�l�ug�꺄 X�I`(4�ޢ�_<��#XKۚBS��'���_y�0�_ƄSi�{��h]Լ�ZG]̸��WS�yM�-N��yU kk��C��'/0gn�9�e�J���=��S%,E}3�׮�A/C�gWƓ-=�2����੷�"��$�
B7o�����.{�_>\���P��Y�#������,�!�����oՓn�&hP���Y��W�r�ci>�h�p�S 
�2��Ǧ�����V8x-Z%6��{[�(C����,���)��3����%�o~:���+�$�O)�4�G��*��K��Zq� ~�6v�g�L^?iE���
��_j��9[9`��s&Ίg��4li=p�����bׂ���Z�V��� �ۆg��gjɊ�ٖ��(��1���Y3�_k��Y���#��b2��#����Wh��E�\���c�-�7�備#�>�����v]��(�^ZF{��_G�d��#M'�v�][�s3���-nםkL�v�J���-��?���Bx�ye~U��mw��A5�,Y�ɝ�~���:�S����{a���{����V�("�3 ����]�ߎ�ʕ\�bE�*�����A��)n�Ѿ��3x�3*1��˪�2�S�Z|Ί�V9�㘡^��RHY$s�Y����0#f�ſ0d���5O`�7Ac��8$>ۣ��ł�c�����C=[Y1{�҅n����\�|�II����b�������C��e��Lh����>6�З0�ۯ%�8{kX���*�EAa�[�6�Y*�H׫�l�hs�"twˑvm��3os�pM{l?��d�i�T���]I��q�n���/^���"{ꙴR����]c=�|O|O+�L_L��ws���Y�g@1��V���tR�z�xO����r�(���?�9���;>-p�*'�[c�y� wUޫ.d1Zt�vѤ�b�F'о���Ľ��,���"�p&�u��͚����9u:0z}b�^����RF��]�r���!���4�w���ڕϙJ��n%X��d\6I�p`&p#Cs� TG��/~��0�|���V~}
�S,-U�[?�ǀ�7'�����'�
�H�D����5kh��\e��~$=jz?B�RȂ���:3�qi sd­���s����AL���@��y#��Z�� ��B�c��γ08�&�/}zHMJ���4�o�H��yDB"4����Q�Ɏ�@��� �d�{���77�'K��UV���Z?-x��(Ԍ�|���o��r39e���Dϙg��3?plIkk�TX�f9�>���Uӷ?˹�E{���Y�)�DvV���˰�7"�?��<r��P�W��;�B�1�V�_G!�Uj��o5p��g&^�eDB6����h34�d�ՊA�|���%Ǻ�����U�ʺL
�ݝ#	�[�D��q�J�B|Ȝ՚�3���T�?])5�c�l��ℝ'D�50�|Lߛ�#?8\�^$��%U�}#�*�*!��o:A���W�}S��(+������%8�����T�yu�.�0��-����~Q�bh`��M�1xA.��щ])Wu|g/oP^b�5 	��+=�jݓy�3�U���)�agd"���]��k�
�W�*g3�t�m��~T&�Tܗ�V��w��3�jw�����]�Dщ��_���@<bKŃ�[�y(�Y���oɯQ��Gͦ|a�=��y}'���"�}�s��=�>GS�u�T�k�m�Y7{�*�)�S���-ʀ�5�pmCc�]|u~�M��*��ׁ��0���9��uU�?���U���ĥ֑�Δ>�p��iaS�k��g��3���&E�d��[Ϻ
3��Yr��'�Edv����O|��]��TE<�"�!�I]��b�T�����xχ�����ݴ��v%@Jl�*��;?ۥ�n�[��-���3'��2����tk9��^}}���f|���:��]�Aء]��_�%���1��X�<P�댐L�ɨc�M�R\&%�cC^����M��xw��2|�!cPr�,���)��P����r)�=�&P:�������K��B��/ӵ�(��=�v�6T}�g��%��V<?��b�<ٽ4�BW�G�r�)��Gs ��80IX�1�~j�({ԮJ��<��v�N��9���N�T{;֟�
���Ts��ٹk�mum��#8}��=�詖����Đ�Xn[��������lm�A��
WR��i)�FS����8���2tt���Y�3j���j��Y�િ+�v�H���1��	E{ΰ��q^>������[���u�(�
�Y�9(fZo�Ж��"w5������PK�'/�2"  �"  PK  ў,J               136.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=Ç_��0ui,���oMiӳx�޴[5ӭ�WO����=1t���DQ���m3u���2�b�ܞ��$��g?�c�-��n��~}"���{���M�;ؿ�{���|��Ǔg	��T/�*��J%,��NN����^H��p=B�e��(��+M[/e5�{o��Ū�K~��k;�ͼ됖���ʑeQ���:�45��V��B�w�%��ݏ�?�S�.9v�z�[��M�~��o�s�����Z�ϓ���Լέ�����6��=5w��]K�L�=x.�C�����:����&:�ZW=�����*̰�Kf^{mmRsXƣ~.������ct濖~�o{�Ӭj�H�����q׷�X��R&u�y��w�m�u���[�3������;��_Gow<Ӥ���օy]�U4u1�¯J�o�[���S�O-���Q�U���4���`�����ɁzJ�t���)2��q]�-�~����!D��2;�s+�W�z��<_η������GfUݼ�i���^�L����>��;�γI7���VYԥ9���%q�W�v�p��ϢM+�m�-���?��G@����ηݱ������	E�2���)}	�؀'��~T�;���q͔[{��:������u�G�G���[�p��<N���{�����J�L�����g?7�~���Uu�*	�����Z���ɫSX':�U�}=�j�ٕw������xr���NW� |��>��ޱ��A4U�~��3y�'ȯ����&FzM��MOJαcj���ha��_�#�����)�g�\�uwו>/?sv���w�g'���(�8���Ӳwb�̙b�����Y;��_�U��.h��$��Qa�����i���&\�[�+��X0��J���&��P�~'��[7�t���O�-y��v��I����Y^|�6w_dʡ��_Ww8��%�;X�:̝��t7e^V��:�`Mz�پ�vf>���?jK��^�(�����en���qu�_�����S/�U������o PK}�D��  �  PK  ў,J               136.vec���Q�����ݝcw����
�`��؊�`�
�`+����x]rY�wÉȲ��rQ�<e)Gy*�T���L�R��ԠfJQˮ�^��ԣ>hH#�|4�"���hNZҊִ�m�h�E{��Dg�Еntw���=�bzћ>����
10�� }0C�0�3���JY����e��D&1�)6S�4�3���b6s��Jc��|}Y�b���e,�Y!W��լa-�X�6���la+���v����a/��ρ,�!s���8'8���S�4g8�9�s��\�J㲼�U�q������]�Q�}�G<�I�O�3�󂗼�5o����x�>�)��s����?��&����wJ� PK��FO\  �  PK  ў,J               137.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=Ç_��0ui,���guO���xx���v��wm/WS￵zݍ���3��ɳk��$T��*�8��墯L��vI�k+�F����#k2sN%�9�������ϯ�8��L�����K��J�9:�g�ui�������^�����h&��pN;�ԋ�J*�yr[��1{�u]|�1k�SNo	tT$�+v��&)w?cbj��xǟ������>�wſ�B7,�EK|{�����*�.����x��%x��r->��q�����{oT�a��w���-�M=zG��u�;ɟD���Xԕĥ����[�H�0K�U�)5Kj�=x�������Ef[��g R�,�t��v�~Æ��m[/lw	ta����[+�"9zf��w�6��0k|W۷����nɷW埝p�`i���-��]F4K��U�@VX6�s}+q1F�>��\g£��*{���)a��2M��_V�!�����Mt'VM�HD$Е.�S�����|�&��<��%\�T�Q����ϱ��]N��X���7hO��S��;I�Hܢ.-o|���6����+�6�-��P"�T���ڒ8�Y�����$M`�����2����}s\ʭVK�gk�p������u����AMvs���Z�#듿A��+��+�}�l���z�gȼÞpF�Ӂdu����&�nl���u&	5�%����Yo�h�/t�5�>�is�9c�����haYɗ�<6ى��{j�X��O��o������1l�����R�ʶK��o��Zw�+�忶��Ω�M�[�]�P��|�����_��얖��Jpo�ik��֗u�]�:��QisV�{��.56Jʳ���� 9q�ԛ�s妉�e����ɳ��N�OfV���ݮ"A���S;/�F<���m�c�������~���e���&�}����_��z���K-��uiLL��o PKh��F~  �  PK  ў,J               137.vec�e˔A����U�������[�[�[�l�l�����%��90��4Y�O�J��4e(K9���De�P�jTO)j���kQ�:ԥ�i@Ô�FYDc�	MiFsZВV�Nm��h���=�H':Ӆ��ot�^w�=�Eo�З~�O���c�>��a(��F�,Fٍ��0�q�g��d�)r*Ә�f2���IŘk7O�����,a)�l���d�Y�Zֱ�ld���V��=����]�f{��~���8��r���dV�S�4g8�9�s��\��,�p�k\�7��m�p�{����G�1OxZ(�3���t�J��oݿ����G>�9��K����}+������7R�PK#L+�b  �  PK  ў,J               138.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=Ç_��0ui,��yk�>�oV,c���?�ԡI#�^����[�/�}S�����3օ�/�J
ֻ�*��*�����-�]ʱ"�ëᮇ��U���3��Z��պ��.�%TRw�ϛz��ױ_W�|�f�8-ԡɥw��S�?��Ͽs�\J�<W��~Ў�5�(
V|���7��9�x�_=uS\���ui���2�¥UO�g��2LQޡ�Y��тO����Ͼx��ga��d�����z<�]�7���^,�J��XԀ[�-:ű�Y�-�~6����vw��{�7{e�DM^�3�</'�ތ�uLQω�w.E��)�	�!|�TM��o�P�[�M�m�N��Ie_-�]?f�&��:Fm�d���1�o�K���tShޒ)�������g�	rUn�;�v���J;gw�o�;���y���j�w��.�]~��#\�~�߬iG�;�b�!B�m>Vy�[I�i����E������Z{�j�kI蒘����J�5���S��ȵ#��k7l�_�k���P���ІRה+jnF��l7io��h���n��k��8"7#���pɕ�[����2���{SmOM�u	0Xԥ��3�3Z�Oq���)�
V��L~��ך�uv����ݲ�V������7O|w�m��w�E/\o�35��̊�hy�/�Vճs5���g�3W�r�����,s�폃}��k,��Ft^������&��Y���hrش���4s�0�1�:�JU��m��d��i�yW���zT�����q���ظ6�?��~���aa/i�����	%Mk}ᵇ3��Y=�]���/�Ҿ�@��C����G3
���|J�w[��ʟs�4���bNJp��4`l�JE��o PK��s�  *  PK  ў,J               138.vec�e�VQ�����������݊�`��؊��
�`�b�z�9.�,����\ΉȲ��PH	-'KR�ҔI�Q֮�^�
T���BU����j�5�Em�P�zԧA*��Y�Fzc�Дf4�-i�"Zgm����=�H':�%E׬8����AOzћ>��_�G�,�b0C�0�3"e1�n�>�1�e��D&���vS��Lc:3��,f3'���v���,`!�X����f�\�JV��5�e���F6��-le۳��!w����a/�������9�Q�q��t���i�p�s�����ey��\�:7��ݒ����|��}���#��'<���|�^�׼��w�=��'>�\|�����}+���H���7R�PK"��!o  �  PK  ў,J               139.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=Ç_��0ui,��y�&�y��ݿ+��u����s?I�]��qB�9�%W�3E���ݡ�����u~�T����x��0����^M��۳Ӡ���7f�������z�u|���Ln���t<g������c����b/�q���N��2)o%N޲=�V�.���+q�@�$O���$�O��l+e�;��e���`BZ��*�������g��)�w=9�����_ο��_�o��ӷ]~�������I�3��9ϔ�R&u��.�E3���#�Zټ�L���:/�і�,g%�ߑ�;o�G�K3��yN��*o=�)#�����0��[E߻gއ���I�5��=M{[�{�7�>l�r���ǂn���Z��=y���+yu5_y�@���o�ˬ����ўi����uC���/V���_���#�ee}�,�<���a]⾏���v��_tUe	t��e�{�~6u�Z9��7k���k��M�� ��h`.�g����[&_��l��������g��(�� �m��+a�����P	�_����zu��S;K��n���#�s���bˎDnC�)����r~���M$ЕΪX�N�lٳ�蒜Ǚǌ��jϱ��>�b��Jຫ�
�^GVE_-1,��,qRsO���x��?�g���bO�8���V�%�J�,��^o�#��������\��k�*fQ���Ƣ.\xv���i[���=5k��=i��ZG:jo����d��R�=�(�ݯ/^q��~��]fs~Q{�����U�t�Ι����>Oݔ�n�ui,1 �ˀ3o�裳+���[�>�|�j;�5e�/���x�������ZD_���ۣ><�h�]1`���j��7PK�_?  /  PK  ў,J               139.vec��Q�o�{������gww��-�b+�b+؂-؊�?��%�bo��p`ND���'G�Q����tʢ�]Y��@E*Q�*TM)��U�kP�ZԦu�G}�k�E4�ј&4��iA��*+��z�Ҏ�t�#��~G��0����Nzҋ���o�G��(��(f ���2���ۍ�G2�ьa,�τ���v���La*Ә�f2��f����2��,`!�X���r�Y�JV��5�e���F6��-l�r�Mng;��n���}6��r���(�8�?��'9�i�p�sn�yy!��%.s��\��y�[���⎼�=��<�q>O�S������#���|�c*�O�⳻��o>�����~�+�PKu;6jl  �  PK  ў,J               140.i��eX����n�n��n\�f�T��a))�I��.A�[bAZ���]���ύ7�Ž�{^�<�9��3��<-<�HTUh�  ڿxZ�p����0q���qqq��		��	�Ȟ��Q3��Q��2��bgd�a�������b`��z%($�K�pqq	�	(		)�h����� �A{��1�Iр�hO} ���D�o���Ё�X�8�x���H �h@ :�5��A�I��/��L��ٕ\ ���"[��B��_VAs�P\��/(���^�spr		����K��+(*)�����C���V�6���=<��}|���?EDFE�$%IIMK��,(,*.)-+��������������`phxdzfv1��{����������������������� @����#�?.t ���н��@���ďE&��m���Y �\�_��EP�/���/��B������d�w`��_d��s-�h��$� g��	����e'z����13s2�t>͊%��Ȧj��p��e곟��>8n,�I�
-�V�x�r ����0$g��S�ԃ���\Q5�2�ҕ���ɓ��B1�X�M�' ���M���9D�r�Ç��'6��.D����\���5%t�D��!�}��vim^$�o�;*~�+�a�}h|h��2����̆؞��\7a�"ε�/���������c?D��\�藫u����%RGܳ��iX|Pa�3������g�E��P����F�����2LY3ґ����}�ú�8t��A��V�fml�L�)�\�ݖ� �����QK�B����I:�۵'=XF�/����Y���N[�,�{D�� ��<gDg�y��qn���k5 �v����Lr-�(PVl�fko�_%��n��xV�:&�n=�zsw�!�B'~r��9�[s�zq��tF�:￿"�w�ڦ��	;�R}�-.���Kt#t��iUyz��~�uà}���U�.!��h7;��ᨬOo�2*��ݾ{���Q%c�q�ې���e��S�
��ʥ�S��d��\�>�n(��C=ܽ��δއ�Z��$�W+���]�F��
����j�/3�i̻UI+x�'��%fd��E�Q�j�p����p�539X��Z	B�t�kԈ�~��YM�/ܩQ�>5D�W�Q�V,?ת��*��OX��k}de/�noLë��Cr�ZS+�FE:��`'�2>��<�~^��N5���^
�����%���`��4X�)k`�qɱD8��w1�q�7Z�XN	��?����8�(��7�`���%�&�+�ƚa��w��xͻ��|㱸�YW��6�x�E;���ĥP��z��b�?�g��ߔ��)���{.O���jHT�ςu�����ɵ�:�e�A���3p40���
�Iw�(bo-o?�8��Ն�@��ο![r���UC��J�`����㊿�n+�(���t� %�Ĩ��>_y��6�j��7�x�(a�%��XA<>��C�3趟_8�ą�H�����E�Ls4����A�\�T��k��e�PYImRސ��OZ�p�s���o~�AX �~3�zg��LX#elǳ
Ȑ��o�[����~l��;Sm?h�Yx���hj@Y7̺�/��^��YNS�M�ݖ�Q��^�J�Ҙ�7�F4�~��܅@K�� �4���̤�y�e�p���,i���f���#���b ?�E2�7���uV�rU������P�Ѹ�a���0k&�b�'��I��^��Dg�d�Ϋ��g ��0	��N5U���*���U����31k�=[7`g�*8W_?������X�p��@b�ϒ̎}Q<K�m�o����Kڲç�m���A���{~������2��Q�M���	���ư9��k��-W�oq�o��<V䴹P{���dݸa�"��F�ըn�"�hx�%f	�ӓ� E�ə2z�sU�I����T���ª��с��7v�W��0�r�D�;�d,�p˃+<JB��޾�w.^��x�׾�������̼��a�N�Ϣ��oL�8G�՞9\@? sh��" ?�w���Y��Z�i�R	џ�-=]�#�&þެ牖��"�l�Xr9�+��q�A��.�_52=[`4|;7u[�3�4�����45����Y�<�^#Wb�ӤK�:"�BkZ�o��>pي-���γ�u]�G��Tl��O�j�c� ��VE5�63q��gB�H�����$}����x�{q7��g������;SzU�,&���l�{'?v�/i� ����*(���4�ɟM�����t���p�e���{g .�Ꞝ��R�b�Ey}�\� I��D�����-h:b��h	=�ɈT����%�Y��Q�]�h��Q�K�bH���-�ai�V�"Mx�b�v�C�m�̏u1�ɍ�]Y��'ߺiJ?�j��qZ3/舼�=x���H�1O�%��{G�3.���	A}.����>j/T�	�k�LޚWu�{��-�^� d��e�Z@�wmX���M����
��0
��ۭJ�dGVd��>#�@<���D���7è�Jx_�D�9�pc>*�������U}���r�� vU~���G5���c�g'��1؄�!�UP$��_��ԡEfI�}���P�ְ��fii�ϻ2�+m�"��D��F�����_�rK�(��J�>u���6!;���D��n�;D�kt����J�>�r0��h&>��-o�I,���z�i�0a�q�+�� �E⢟ !^Gۊj���> ��+�ҋ����e�cE�4�t��#��e�M�z���WS�a4s�i��h!����z,:��&�B~�0�X7µo��Y�	�g6� �܊*�V?Xa0��NŃiYm9 ���p��m������T(��Q���l�E�8�����`���ݝC'���;����!�BF����i���z}7��fQE�#�L%Կ����~�,XP1�"y���9�_`����$xB� f+d��@� ����ib�&
}
�V/�ET�oZ2�\H>��.6x`/`�$X���x�k�'�?0BK�;� ve��Ѻ���(���aX.'#�u��ڇP�BB�#��Ÿ	�ȏ|@���7�7�ƶ�>RCK���R�A�j�R�՝��S������|�~�9\�S8�/ߎ?D��w�����r��X���QV���	�i�f��M�X�?���5���%��T��K Pa4�/���[��'�|� ��I/:ĉ�d*ܝO��tm�0�9.m�^������O���i�m{�͕'��$���$��^c^��%�,�>�)��µlHW����h�z��2��½���FE����$S��<h�QM㆛í�e��1/��D���ڡK��t�8\Ԇg�{�����O��B
v�Ip\��C����Ā�!j7MO!#6�&C芷��k�l�<�}��C�ʁ`nPI9}�mN�x=];���_@����+��R'�y�4P��q����#<���p{���=�a��Ui��v�{O�ݓc3��Z����BX/����`����Y������~֔�w�[-D���X���lX�pB<���3�E������o>E��,�h,�@�
s;]��sw���R݉u�)Z��Z���s���TZ��|�	�������y%�A LL�tD!�@}$��p�O��,�/�r�H����*����e�5��)P����:M/��U�G��=}�Z+�-����6�W�r�UQi���=�=�-�[�7�c�wN��2'�aAa�aڋ��J٣,�=,,�,@`U2�([�����)�����T@h�zI�T��yU����4��$H��Y�"�p��}�1�q�&n+�jL#$	+v�h|�4�XOj�m^V9��f`.[b���t��5L�E],k�0N�ܑ�%�e�� ���y�����J��J7���	t>����pv�{��g�$Zv�Z��@��/��C-{��1��	 �V? �2u7��up�ߦ�kUvPV�tiJ��Z��-1L4yD8�i1��I�z뵎=�D
1yZ/@����݃������wΥ����J�s�$��"E�up�[B7�%S�B�j]KuO���a$
D���J��uO}����Ex��K9�G�(��{e��u|���c�x���bs��>;�G�#��t)�5)xJ2�d�(Q������y�h.��A�8(�.E�leU�����v�Jޏ�9��[n��!�����d�a��1R�&h�Y�x5��č�P�7I{���;6k�ΩM)�-znCI���������G�%�R�L���%�o��)��S��WU�Q��9�� ��r|�����+��5�'F!�wAya�C)�?:�W?3-��Qb_�@^wJ�`(v�zu�7!�||7 �߽(��P�.W
B=$��w�Mi�.e�T{��RF��.��p�^�p�HT�罹�����F9�-�ڂ>�R᫄z���}\�� ��e<HuX�3�ΔX���q����"�!w߰�,�(�i�X�2�q���H�r��}��G�\�:) UH�b��M�x��X>�n��_���FYj��R{g�ޙ�|~�&��5��͂�Ư�G��"��e%��f��5��9�^k%Qp@d#	~=E?|T�|�ĕ�9����n5�)�Ia`�7��U���˝}��-�tk+�?�C��	ª�>�8n��%Vf#�bSc���*��#�?������ƫMW}8�[v�.��E�w�o�^L��~8��
x��O�j� �@�o	���I��B�"���(��)Q'��+��o�����;����1��A�S/��<ƒ��S?Ij�O����f�6<�����ơ��I'
Vdsv�Ć�e��r�&a�M��`��gf�Q^m�� �[D�-�3��}�ſSM��kJY4�J�ޘ^���+ǒ`(s���X{/&~9�k�����1�?W��C�8�S�8��b��&Hڛ���!�ӅE��H8�^�&2�l��:v�c��Gz_-ZW85^�ONN�h��w�3����!�֊v�JZ��i�?/��T�����򍕗��@�:�w��
?;��7�|A�R$���{�[{�Y�͘s�t�!^(�4��\�)[eY[o�0#^��_�r��sy;w�b���@��W��,�Ǡ	�fwF�G'�| {�!$�Ij���J�(�h5��k�nzb.����A�p���'�UpQ������C��"���#��I�e�v��`ʓu�9�������Dq�Y��j��n��ce�%Ҿu�1��智�p�"��(�"��B�"
0���Y���򃮇�D.�����F�.�/�ok� �����S[A_�~�}|���ܙ��S�`�
��Te!���W	*��)�w�~���`�\�d��\�g�J<�����lz}��X$9�>�έl��b�i'y^�
L��#��1�Sb\gd�,	\-�����v�/��;�:6bL�5��*�-9��r�MB{��V�x���в��UQFճ�3�qM�@\c�p�����&̣�\'�}����&�;	��w ���WdHowO5!�'��
�B�vCH��_!�����zFb4� ղ������R���0e���-�����qs|@٢z�B�Q1�C	�N)0Pm%FIE�t��E�f������`x�� r��rmx��a���AM$Bp��s���>���FR�7w�Zo�Bn3Ko6!�b���0A���pa=b���r}U�N@aްÿYy�
�����t3>�8ؒ�N1�
�+��T�AW��V|OQ�ɂ���H)E�f��&K�b��UiR�>wx����A�Tl�R0t�W��6n�=��"S���实%�D�2ȷ�w�d�9����xO�b�Ѧ�E�^Z,���~Eg�#㨇fzݶ2��\J]<�b�>�9Y��� �%��t�BK��]�gG����M�b�QF_OI3�w���>�5��絪1NmQ�+��DW��-n�
���E��&@�)Q)��ퟺh�˥��&��-ng��R�]�<��R# �x��A& ��y7�yA���ktn67���M�t?>� A{�� H�/rcפ,F!�6�G����Kld��8��oӃ�G�.sjBɱv���ؾ���a���K_jJWt�|B�z�(�S#�4�+�޼��A(nO��;IB�*�K���钨����V�NU�e�1uK��e���'}5�S���mЗ%�^���L��ðh:�D�S�������v�,���4���sC��0#��0(��>3�KA[��An\ ��,D��g�oJ����k|W �H�$M��Ο��1enGқ�nh����#S؜G��w��~�[(B<�\2ƕ��|?+ML� ƽ�6��B&���4��Y�����D;�xsK)&��W3'��b�d�U�㋃�*!G�7�sBB@�v��}Ԓl<�t��pP��u��s��k�4�M۳ߌ����P�)��*9���8)S�g�b$�Ç?lW���\V��%���i?h�E���Pί�잯����nc$n���YCd��;�R_����.��bD��X�BNPw<S��dz_@�A Q=��͍�$7�7\�8���,�V'��y���	�:�H��7�}Aa�n��jH�#r�",$�>V�����������������Ku�c:V� O�'Y>*(�V_}AХԤ�b��ɸ
�J�-V�W1�t��j�W���vyJ��	�=���'���I3c%_�h�T�~E��r: �����O<�3I�9CfZ��a����r�[��w��'��ym��9��)�{󶈇�C�ی���u�
QS���b�EEvv ��,�wb� ��oY�N�uB���Y�O����t��mT�T{*ͥb�X�j��}y]F=U�(����[
�3Y;���_���k�.Z\�i,�8���Y������:�#U�E.���ٮ��^p$GV"��P�y����*����Ge��Ō��7yr�ZR�-+ڭ(r�!�V/�;{�s��n�ɩK��9Y,�_N��2[UdP�~���G�E)n�`3��ˏ)�g�H�+���\	�f���%
�End##	Q����t�`[�NQ~�m A�}F���IZ�	�ԑ9�����%��w�I�D\�����~��2p��O�����MFH����́�6}ql�p�6��~�Smр(���`��ʠ�&�u4M�{�Խ%%�a�I&�ۂ�V4��.k��)Qk�_`�]�	2�1�B��k��r�!C ϳ�P,��=r̖�MV�9* ΞV-��L�u���j������Rw��FK$�zv7+�+`�"�]E�x�w��Ź�Y��8;;��Z��U�o�rN�j��I��H�٤nf���:mrr�,j�7_�l.���	]2>~�W �=Ŋ��y�`M�T�s�s�t�1ɋ	�FiL2.8�V�j|.�b5��أ)�!�Bw�Ӈ<),�5��ˬE�W3�6^E������f9u���F⑔c�F�*��3�[N-���X���d�0f�F\� ��>�����x|��FϩF|�~��0]G]9��ߐ�롱�s5�K�>h�}��qH7�Ԋ\F/�:��OW�Q�0�2W�9�ڨ[�`J��ĎY�Z��Uwv�OqN�ڲ8��xzx~�a�d
�.�2LW~,}�p^�~2y���Y\�M�Z���@�'��">W�o�?m�J�s�o��BÑg��YTJ��8Efb��}^b�'�B-E��!_�+��8�]W���?���Q�V�Jp����^���2��b��s��1ZQӇ���OBܩ&RNƻ/���Wӻ�n��T;�sq_ 5Q�]8͌�)��c�#�㎷޷�ۭW�l\+G�ֈW9�љ:�!	_مӠП���6�۳�_�D��9zC��"R.8K�RHT=�>J�7�i�6��e�.��S��-%�2���AHUk�����3��+����S|ij�V���Q���B�7�a:	:�5Ȋ1@P,Y=�M���0;+��U��E_��UFF�\�����F1���<ދѥ$&�-j��M�*�,H_ꡬ�E��	��cu뚩�$ 6�B�ͩ�(9U�-]7>.�(��i=Y���j㯣�rk<4l�ti���
�tG����_	�'��=�7Y����?d!�"���W+�$����X�����u�[�M0I�t{�}}O�?n�(��\�a@��8<�M�$�t��#��ɀ�mzy�,������($=|��X�9k�"��j�a����F�~"c�}�lѪ�- �2�әM����߃��♯/*��i�<�T��a�#埚���UT󲐜�l��o19P_���$-�����7�u����a�(K]6m�=������YR�V_�*��Z�$�'�;�u*lQG�j�-y�2}]�5��'(��8l9!G1�	l-j�їgE�,0�tQ��U���ʅ��2�z-!3�c���޴2�>�i��2�IB܈5ߢ�r����+�	���#����i]����lj�w���1����~�PK�r�!  ;"  PK  ў,J               141.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=Ç_��0ui,��f���g����%mgg��i�5�/���� ��h�����~+n��;e�K�>���B��<).	tTt	`�#f������[�ѯ���/�}5y��r�0�^�2����������*�3p=�8hj�9�l{F�~ނy����<��z"��R%�}aO��i�!QAO��'�s�����ؙ�����҅��z,Xԥ��3����x��8�/��:�*b��ܱ�u�x��bkNN���y��<��1&�_K����׸��S'��H����Q��.s����e���s�|a��z������-M�[�ªKc��Ƣ.\�����Bw�OԜ���v����v�t�;|owl^���Ni]�&��V>^y�����������lu	��)��V^{�vٕ��ƹ�">���.y-����b�R�.MX,�R���ߪ�W���Wy'�Ui,�q�@:��?VuG@��[����9���B�|O[��ȭY��z*;]�VjX~��iތ�N����AY����}���$1�٧�����)�yR��颗+f]�澶�8?`�����b�}�uU�3z�_����@W<�q���-���K��N2��.��z�c����s��z4�^s���W�q/�qy�;�]sC�V����i�n�������|{r����~_/%-������?���m��O���</��u���7������#o��ky*sͼ�N�P�f�u�6��(��ʾ�wgN�,��Ͷz���������ɧ'L>��|��ϑ[>Z��L�}']-(�]wZ�K�]�_ֱ���bjr���<��$�5�D��������}���>�zg�-#�yi���ҙY7{�\����Ďo&7�,��Xb@(�m����f����N��*|vw2��|?�V�}��V�wD�yy��w��>��c��;�ǵ�ģ�_�3����*�A���o PK�yVi  s  PK  ў,J               141.vec�e��A��=�cwww뵻����l�[�[A�؊�����2.{�̗��,��'G��S�2��\ʢ�]�"��L�R���H5�j鵩C]�Q�4���gM��4�9-hI+Z��}m�����@G:љ.t�[*D�,�zzҋ���/��o7�n�>��a(��Fڌ���X�1�	LdR��d�)�T�1��d�����\�y�|��E,f	KY�rV��U�fkY�z6��Mlf[ٖ�b���Nv��=�e�mȃ�0G8�1�s�����8��r��\�b�7.��\�*׸�nr���)�(�w��}�G<.�|�3���/��T��k�ؼ��x����S���H�%������?����PK�vL�g  �  PK  ў,J               142.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=Ç_��0ui,���[�D�+��A��'i~{cs��������[6DE��������Gԋ��m����e�fͳ�suiuri,j�'6�j�t�cr�������w�l?e;�|�Wu=xE��S5�3��q��v
�%ͼ��ۢ��;9S=�'*��?���l��>F���~O��Of�M�Ƿ�>���.�sW�Z�H��.�E]����|�>.�ؤ&>�2���t{���g�y��Y,	|ְ���?�׃'�"�G�H�_�Vq�E,_^,H��N����}��^�[g�|[~Y���s��'�m��1����R��0�@W����2AǕ���<-�Y��zx���Vv�]���j�K�+�q^�~����I������`xC��*�E3XE�aY��oWL�t�a��\�M�?�K��֯\����a��*�6M��)jG����^��wڊ�$��0��쾏�9���і2��ݺ���ӟn�/��r�ge���ٝ5�BY�;^�z�n��.���\��Ѻ��Ţ.nB�Ċ_`��33�}1�
����L:nz�ǺsҺ��g�]y0og@���=u[�����w	�&�ʀgULzs7���	ݮ�>�����ױ��Z�������t]���^�Tv���{��z�I�ӻIA���Ӫ'�a�+��s�W?��[�����e�a٤B�����6����]�O_���3��qQ�ץ�e�;ME�#���w����u���,�j��k�nޏ͏����t9�����[C�����^��bjWu�D?�Cy2���V���=m�Z۳k{�X�~�+ۛ+Y�Qs�����w���N�y���e�����v���t�<9�zǟ���y$Z�S�>(����ю �'��m�Roi,�p�@��w�Ƚ�]���r2Ş/8\��S�:�b�罽U�ͧ��
�~k=�n�Β��qs��?_�����V��"Ax�-��	 PK~���x  z  PK  ў,J               142.vec�U��Q��]ϱ����[����l�[�[�l�Vl�QG�v�f0��|Z;"���+�9��)��(kWN/O*R��T�*�R.����kR��ԡ.��O��0�h�7�	MiFsZВVv��\���Ҏ�t�#��L�T��Y>����AOzћ>���]��@1�!e�a3R�b4c�8�3��n2�n�>��Lc:3��,f�?1�n�>��,`!�X�����`%�X�ֲ��l`#����fE�Mng;��n���}�f�<�Aq�#��mNȓ��4g8�9�s!��%.s��\�:7��-n�㎼�=��<�q�O�S���LE�J���[���|�#�R>>G�/)��T�����'����?PK�H�.c  �  PK  ў,J               143.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=Ç_��0ui,��v7�C��>j���~×��&��>�~sZx�M�Y�SXo�{�@ �����;O��0���ѯ�EB���I.�E���J��%Ź���+�3�Ӟ~����uW���\�g�,�HV(��=A������흹��VVK)����Z������=�;P}aO�X�_���JH�_+,�g���#o��}s�LN����D]p�R����V�2VSah�i���(�=�}콽�ܯ޼Ԛzf��'˴���L��f�e�s�C��$Y�g�V�d<ϩ�v�������'¾�=�fk�7��y�Oq���y7W�=~aץ�ZEcQ.���u��.�R�rir��[��6����O���	��Æ'�z,ìy��R�Ƽ�E]��8c���d����]�0و����Wſ��*9���u���jk��ג�:m�C��+�l)Wۃϝ ��&>[F|���$?�����v��]"{�lI�B�F㟛>X���JǺ���E/
ԩ|���jwm	t`Ń�g��bl<�Q�ټ=��DOm�g��&�G0+�d��['��ٓ���m�N{��U$d����S��o9�����򻛽O�U��u����w��R���S�������9.��w�8����l��;�&mS�6�nEDV9��=���w>�׸x����2�=�F�s�����K{�X�gv�Ϣ�����U$  _��v��Z�@/>9Y}or���e}���ov�ٻ,��j�ѤPa�+&�WwǪ^Urg/W�8G�����������6��!�ߎg�؝�xN+�'3�==%Е�Pֳ�->����������e�c�d,M�W�8s��F��}F��~��2I;�ʘ�my�afY���E]x0�.A�f֪�	��*�|@��u\����E_�������)s��t-o�4���x���ԓ_�3���RW|����� PKܧDY  a  PK  ў,J               143.vec�e�Q�w�����[�����`��؊��
�`+�b�:^��k��/��DdY�r��$yJQ�2�MY��+�W�"��L�R��)5�j굨M�R��4�a�h�E4֛Дf4�-iEk�6Y>���hO:҉�t�k*D7��zzҋ���/��o7�n�>�"3��c8#lF�Q�fc�x&0љL���Oa*Ә�f2���O̱���c��^ ���,a)�X�
V��լa-�X�6���lak��mr;;��.v����s7��r���(�8nsB���9�Y�q�Yq\�����r���-n�㎼�=�{�@>���x"����e��+��76o�;��|�}�_R���o|ӿ���wJ� PK�k��i  �  PK  ў,J               144.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=Ç_��0ui,����5������]��.�ctBb���Q�c7oi��u���c�3�[�)v3�&͹u�آ.�I"����y��>��I�,a�ûhg��eV�<.w����l��!��g�L��_W�,+��np]��e���ڊg���܂M�����b/���S�k�3���/�<g,hM� P<�s����,�E��"��8�l�V����+�"�b��9�N����^�����1{�rN�T;����Tt����#��o�G�H/^q�r_�	%}fY6��E������{�ڹC}����YG'���<�gT��c.��%�5R�U$�fO\���H��^B�qՎuB1��]�L_G$_�t����g�vu�#v<�喛,��^tU$ЇPb�[|��ٯɋ�lY��}p���S�����[p]|��b��)Lүg=������G�nVMt9F(���]�O�z�F,�<W�b�ރ�M��ϖH�����iI����yAA����5�s,���舾��U$HGcQ>|��z�K)O���,�}�ul{�J�Un�5��wD�o�g�t#wY�-7u�m�/�6�[K��^�ʹ$~��m��È�E������I�����K �x��]m���p^���L��(L�`ە/�^��������l�?C꽞m�n���r���y�˓���:23��B�}���Y�L��f�R9�����j{�]2�6Xíd�f�#���:.���{��$V��{OC�W:a�=�\ѯ���]q�aMԍ�y�>�����m���e��܊)Uy�U�HEF<���8ݦ�?���f6'�;��}���%���ј��=>���2����誈/�@�ɾK��C"�O�+w����a���E�3�4�ӷj~f���O7��!�G!��P�)�EJ���\Tظ/SƳ��I�e�*�/�,��U�
���̫�ɦhO�����}�]��XV��\��R�Ţ.W|.a��7PK#ސ�  �  PK  ў,J               144.vec�e�UQ��̝kwww��]��]`�؊��
����b+���;�}��և���Y��"r���@ŔE%��z�R��Ԡ&������]]��i@Cј&4MͲ��zZҊִ�-�ho�!�EG���BW�ѝ�L���D�M�ҏ�` ���`�!�P�1��d�c3V�c<��$&3��)�4���f2���a.��b��B}�Y�R����d�Y�Zֱ�ld���V����t�.��=�e�9�A����G9�qNp�S�Ί�<�9�s��\�2W��5�s����n�;��^�,J�}�G<�	O�x&�󂗼�u����w6��>��|I��)�����?��o��7�PKf��c  �  PK  ў,J               145.i��UT@Ӧ�!�w��Hpw'Xp\�� �	� �����4�������^��ۗU������U�+Ͽ DjJ�J T  ��<�^�01��X@ ��������������������%3--�8'�����;HFBH�OXD�?��`cc���Q��S
1�2	�?�@��"�����J��F��<`��'��?������	�������B@EACCEG��@G�g�g�c�0	�c��� _BȄ"R��������X�m�#�q(^PRQ���spr����K�$_�VTRVQU�7042615������������>6�C|ZzFfVvNn^qIiYyEeU�צ�ֶ�����C�#�c���K��յ�[ۈ�ݽ����˫�7�w���B���O����q������Å��bt&ALy]����P�BjQc?6��������o�����7��X������\k <4���F Ή�}�U�TlG)�w�1V	&�4����Q��3&T����v�m���0<�U�GK��t]W�ge_-�ξ�Uc�Mٔ|�"os;m����nr\�����)�|��G�ֵ��R���2G�&r�n�|,8G�f��W" p��ei����;U�y��hw�w�N��π����\� >I�΄*|���v~� �ٿ|R�[n��>��AW&��ޤ�I	&����V����������C�7�Pl;������"���͇��e�:!:�_��'۔w5��K��q��N�'��{UCN/�~i�l�R�#�$���Ix�`X�nX���>ũS��M֖� 4u��!�j���Sm���Ͱ)�{eҰ�T��AJ�&��0�Lt��V��W�9`�����R����濥�r�g}�F���[&Fi�1��������t��W�҅	Q讧�Qe���%ed�˱;� �Wg�\��Rd\M��?K<r��,	M�)QK��F����מ�w��λP�9��5����zsH>M>�?S�|�d>s��~��➭+^B�g�G�3L�0sd�����P���Ι ��K�7$nX�n�&1&��j���W��ӫ��-�l��=����C��{Fl�m���U����8��u�yfs� ,��^ǡG��Yq��(������3��������n�>l��20�!�^Z����\R=mXc�%�Xp�M��0� �$v%�����Wzq�WE��rN�����1����d���f	3���mXlk�7�d��v)�Le�7iz��^Y�֑��*-یh4@�v}�'�C{��$/�҆�'"�*��ir���c�	�F,�7z[��ל��o���]m�I���	�dT栾r_��<
~I<�(1�z�~�G-�6��
�Pr4��6�b"�8͟7�v���s *ߨg���sd
��������h8S<����Au<@�4-j��m8涝
���.
'�ܕ}Գ%Hb�c�����]<ߖ�ƙ!� �b��hKq�+�.��f�T�H�&�b�85K��لp�E��	�2�D���7Ӈ�nB�d����6:��~y 2�u����$�.T���l7�̣����e$N	��]��$L�anN�r j��2��}F��m���ޖ��Q�L� K���5;<�Zp��hO\׏�T�P6\̦i�[�:�urM5�i� �qaj��_���liiS0����t��?�j�ɺb�4�뿭���F*�p�4<bȣ���\)��VX[��t ׈eխW���?��D���^��|m�b-�䬁7��o��׆ͅ��5�N\4�+��`֤F*C�_�d�p�c�O,k�`���V���>&M��(�	�+�'���7������)�K�3 V�W��gҜYT`I@e"�������Mm'��FS`k�I���g0��n��d�����!8
g�2]E�Ui�3���&�ѹz����kNk���?$lĕ��9�$�5@��cv1`d#4^�^�t�xj$�7�֞9����s���℮i�KT��|٪\b5L�f�ЮB��>�w�������fqF����Dp9H�
n����$E{�'Ow�=4�(>�nےc�/�٩U+E�?f��%��ծu8���\�6��$am��|zP}�%��v90�wG�!O����e,���hs�x~�C�ߘJ�b�?�N�2�2��c 9T<��V�j����������,��9����J��y�=8&�O�({���U���ϗn�?I<�m�T�|����V����\�xi�{d�ss//EY�P�1�J��t��5^������(?]A��39�Gy�2O� ٭j��,Y��ӑ��k���bT��F��tF����䘧����&���ݲ�d��tҐ�.�w������W!t��U"��4d�Dt�;�b1�'t,�0{X+̟�2��H�6@<tom�o����F��%U�j5�ݼ��5�b��/��R$һ���K`�v�g)YUؿc���w�>vP�A�M��� ;y�>9�3��'E� �DFY�2G�.�-���Q�y��^pN�~� ��Y��s���da�k�)X��@j�<rއ�.�A�A*Q���kq�G�py�R��ֹ��qW��VH�12<���-~�r���rdyL>��'�	U�\����x�#dr<��lç2��ڇ
)�[y��������F]Ɨ>�X�ao��#x�\�ׅ��T�G��B�}�����e�Ӥ#)��$�X�j:�_��[����)�A�^� ����]p�vm�<��I�.�$��`j�b��Nl��,�3 ��6���T� �@ Dy��tX��Q��0Aˬ΅�����9)�qbK���A��޼��{:7Ks^E�y�o�_�6A�t�����[�\}#,2;h�
�x�p�.i���lI���ɏ�5�7�y˻.�N�c�K����G��@�'��ߛj�� n5A�r��5��D"�N^���I�{��
J��N���J�4-��<�(;����N�0-q�Z4�呋����A��tb���?ڇ����q M��e����?yҢ$)Z�1�{�$�&��)�zr.j��Os�%�gƚ�2>��-
��8�����eЙ#9\~fO^���+���$9��g �C�3��mlZ�.C)@�sF��9˫e�S"i��ّ�����1�XƤ�䗥w)O
B�WG����׭&��&0���j�q���io9�T�ga�C���w�,��8�6;s��
߻ocݥ��4u,�����k����ַ:�5L̷q�{�U�ꪡ�`ޥ�z�vυ:�*��k��I�d��~����
�m�ܛY�V#�k�#3Ɛ�,fA-h'ʓ����f)S��Cƌ|��u=T��¸�l�m��ٜ_Yx����`��x�����6�5Y�r�X������X��86i\�p0�|�̴�@���U��QYo4�c/W���+~=��� p���U�j��a�P��
��f
�V�T s�O:�/����y=���2���ń�7Z��`"w-e��g������(3����Dښ��`Z�^��|���d�l��n���Q�*��i�t�*�_�S����3������>֩3�*��Vc讳���}k��y�9	����Q�v����Ǩ��� �I�% ũ4-٦p^�F�+���e$Ϗ�綽Э�#�u~��͗�P0U�=������+r���F�n��@�]7K�0.g?8�ɥ.�qħ�C�3`�Ye��R�dK���|͊���4�T�ޛo𽣖�Y�O��`_��N�pUY��`�_�?lS�\!�T:��9�%�}��\ߌP�2�w
�`���=��/L�HK(�~�-��
����~�Ęjx8��iץř.!kw8��A���m�@�K�!����-�|���u��b,x.��@�mA��/��7�o�F�?T�6q8�(#'z'DʛY=|��_/���_s����BV�����<����`�pc�厉5�a��T� �	z����*٤���	���� ����p�VEO|�ְ��J�,���������5��K�Ų���5W�B�7*T�t�9���{iξh�>R׿�Y}�F��D���7�a�H��@�p$II2��Q\���r��x��l.�#7R�3{�E8��?��ų�<��K�]��x��!;�@or�n�� o�,I�,��f���&U�s�\�d42p�Aaj�
g�.� �B��Er��3�b��d�d��ٍOcG��[:R��*)~]�� kM��%ɐ��w^%:ۨ�EM����9�+�+�&�Z�|�@��0�F�=��Y������Ficp��O�W�R�|�i`�>���X�����D�{�ln�xck���[W�����o��#�[?v�X0%�.�@N��m�:�ż�F�3����`�.�ߥMO��!����{|ڤ�Pc x�<�*FX~Y7uLtb$X_��& ��b<�O�|��pn�U#���g�*O�(�+�|�\��Ũ5\{�� ��Y�EPf��Pc������᎚j3�(����o�x��4��&p�_IO����p:
�%�fQ��K������&)���&�Ν$���xq�u>�N[Z"j�A#nG�����NQi���e0<�d�{��t�TEy�H�^x�	ut-Ķ�;^�7�Y�ˋ1�?����E��!�b��q��2���K��������n�zff�JBoK���Zf��˹Ϣe_����k�\��g�J�93����}�[���;��x{�O*<����(<�������"R�Ӕ�)�;��m�Q��$[q��1���`���`�i���s{ק���7�e����
��IA�d%�}������&��vq��'e^�حA��/��,o�����=̥p^�D<ɞ@�8��|�|M����TŃ\���g�!��J�K���T���t�Q�c���eW�-�U�xsI�5��Pf�?�<դ�K�2��Ȏ*�;����O������t�K����(}_F�(90әlu��Bq%+=E��h��5�%���
�oGd^�u[�j�SM~&��@��H���dW6-5>F��2]��ޑp�a�	P1����ߪ;p��z��d �ҏK�Z�!'xt���/vr~#g��h=��=�\(!1�ث��ug�|�Ik��l�:�exR�׺�o ���idj3�
�]��2[G�J�zC�����GG��]~�̎i�k �DU�hfg&��c�cYp��_�%��{��>�fK�H �	Z��x+�ND���
�w����D/-ug>}��mU���{���]�Έ�Ǒ6�I{&\G*^��E=����fqn�ko6��e���(�;Tߟ�g7�>q�my��9��`�/'��V�!Π@����H=�,G=緡�/��Δ0X_|�T2ڏo0�aw���`c�0�������*@�s��[��C3�=�f��O.��O�۰�R.�=��BN�8�=R���$?9<�l����u��uቯN���rA�_V,��^/z��g{�S�[�R�VF�t������{����G.�b�/7q�޽� ж���l�;3)uu����`���꺪g�Z�I3Rڠ3#�t��\'Y�xg`��` ��I�x�*��־�ډi�L����8N�vYY�����X����h�]{�^A�ީ�*R���>��+�%���D����1�FG-;#h�3�e�vпYv�[=����,��['"���pf�bk���t=!kҶ=��˟w�p����H��h�&�v�h�?��H��W���"?*6���Sl3D����5Ty�?�K��As��<��s��>5~��A�ݻ,���O������m׾����hN|��mIy�_1C�Y�*�l��p���E�n��I'խ��٬y�
g�����s�~�����wޖ�!5�z}�b������������y�kf>GK�%�����#뱣Zm4��C{A����e����!��K������:�}M)Nh�����x]�.fZ�Mو���b�/k��gM��|�!{��iB����C��0����SOc��$�D�F�6 j���Q��ރ��rG��)W(:VI�Rʩ�I{�!3G8�6�I-�v�����Sq/�GY4Z6C��	�&�E/p�l�-:�8��ĭ�yބݫI�n	R
����h� �*�����2c�BD����b�KP'���a����ǄsyY'&;�o鞀�y�{=邥ziD�����)��v�u;쭕+D�����3ʰ�F�D��0?�BF��[4�0��Ks�,���E%��
}K"�ѽ�X�򉓊+bQ"�+��ѿRO9BL4~¬���w����Q�������a��R>�f��H֠��J����/	���T�-T%9kȑYnS��ۡ���������zI��{�k���s�nUa���h2zL�g �NE��B������K����h�`C�ԇ�/k_N!IKj�aw���ݯo7��G������-�<�/N��T�ñ���.�ߊA�{���rڊ���M{�uߞ�>�'����tW�2�J7	�	?`��Ȁ[��!�}�Ɗ	t�`�o��� N�ܖ��ټ�A�t#�%��*�p�YApl�¥�L�uB qEn���&i���au��	 �f�}��pWm/V�����KE�g�������ig�I
���������8l�#�)���{|��}�m��|2ȩ��	�����u����)q�X-���M���H[�_�u���1�uO�N|�X�n_�w�u�ՎG�/>9�~0o*jNlf/k��}Z�S>q�4F���gΦQ�π���5�]���wд[y��X�4�ȃ���
5��Q3���oW�#E�v��{��@�K[A�,%#=�HC�q��gl��>��1P^#5�Z�I��'�ݣ��2Z��Եq귦�ѴO�O���8���PQ)B������֭��r3W�M�eZ�42��4�vI	�.��K>,�m'����'�W/��Cֱ�j0�l�����]A�_��f*T�k�[o%<��c�Q�?��s��Y�>1jDFS�(᣷�*I�=�4M��xY`����c��1��I�x*W�6;_F�j�5EE�<�~�U�V�b�"��+���xԓk��Jz�9��'������8 C���g��^�Yf����G>���/�
��\�L��ۗ���~����Ӑ��/*��π��-�2��Օ�~f�����]K5D�6Y����<�S�y��֔f'u)�E?eے<����lc�ޝ�Z��9 qXlX@	�s{���|)��ߕ߸ע[c������5�^��QdI��"�H��'��{}T��n�..y/l�qq1�`ܨ$�v�a8���r�HsC��\G����c8'��,�O�;�%���r�1��1���<�7f��Dg�\Ǐi�y�IN�� ��y�-D�Kd��3���r�g�'��A�Sњb����l���J�[�|�>������ �J���kG�f!u���nij�ٳi��l)��Y���T�1�{��33B���m��M�����j>L7Sn��y(��g���[�K
��B%�";S�f�v��1�.^υkv&i
�����x�q��ң%�b�"��+%�UD��z�Ь ��D�G�@�6����@��7b��n�b�"��d�3w�{z+P{���;���.fm;:��7�euf��yWd��d������f9ͻ��[�������kLO��}
���;�_TtዱxW�ߋ^�~8��1��s�7423[8��׬l��ӋT�L�-�1o�����=�o���Bd�d�k���'���74ͷQm�,�u��n�銬>�%L����nG�2�Bfz���d�_Y�M M�R<�׮Q��K�+���L�2j��=V-�ߵ��ĥ}�9W
˜6ʏ}m�4��qq8��qt����H-���[���������x�������?o����� 쮟(7�EVur���,	&�o{^�y5f�U4��E�p���_^�+����N��b9�d2��2
���|�T���>Giv`�H_�T��7��E�
�������Y����+"�ٖ�����(C����祐S���y�.k@r��^'��O+�j>�0o&-v��E�Hd���*��&�6��<����_�h�@_T����}[L����8��~3A,j��ʇi`��jW���UOtT�ϔ��p�kff�3Z�S��}� ��VU�b|�n���#�:��"7� ���p�����JTS�fH�`�uȅ3Sh�=��5CeѨ �)&�ݣ��шYE{����]`���,�yC��Ys"a�VYCʌ����9N��lJ��������ϐ���@��Cx����Ѽ���h�9�$�䞕e���9�A�[��2B���,�11�d{�/j��Z���-U�Y�I�TQ��E�wz!��o��N����HO�y�� PK�+&�!  #"  PK  ў,J               146.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=ÇW�&��:�b{p�Z��k�˛7NzR�̸��%?ׂ9)�}f��,:{щ�yuS��G�۽������g+�|�5k6�_�ƨ.�U��"tČ^r\��L�._���N���mWsk�:.J7���ڿB�g�:��_W4�|�s��������s�<O~�a�����3����x��T}���W�P�ݲ��K'���/�t�t�XԵ�KcQ.lu��Ʋ5�u�j�E|�$����ur�_{��{�q�p��3o�`�v��:%���זY�oس�Gx���37�]L�r.\�|��k!�7�L9Vppc0����4�rⷼ�U��麟.n�?��I�?��+�Y{lwi�ڊ���m����zĩ��Mm�5K��Y��FW� |�=���ū)]��$Ծ��zRs�<g֫?�W����8��s�CE�u�n�i?�[��*�Rh���.<�y�G�����:�.��OҞ��:�ӽ�n�}�H�%��{B��'hO��}�]���i�;��4l dr��	w#��9'�4f��_�z�+�f���z)6Kz���F����~/��t��ݹ�K�����'+-oP~�6?�?�sc��Z��n��p��p��S�Z�Eh���f`T�_��Ȣ.�|	s��kKO.n-S`�U���U��[��	��G��V����"9=��f��	��v�=_��l��C�뽓�g�t�ۯ�x��=�&.���&�t���I��T
�ڍ��u��$�㱭��t��;&�<�3�k~@���E]������ �G�W��YZ�g�4�ڲ�*�Wߕn�ٳ&��6�����|���+�0y3��%�<p>�����c��Jk��<�[v�O�����^w8�>T�eᆛy��I$���y�T���Y�Y:�{s�?�mq��4)X6�T�p��t#�=�K�/-PHK�R�0�(�+�x/�2�V�z;��&����n�se�®/���Q�zʜ��)�q�����:._A[i���DىYXӼ;'l�n�R�j�D��Ò+B%'X�����js�-.�&>�b`(cH��7s��gF]K`I���M PK��6i�  �  PK  ў,J               146.vec��a�w�{�����V��.��][�[��l�V,�u��G��s`�TD����9��S�
T�Rʢ�]�*ըNjR���I��kWO�O҈�4�)�RD�,-����5mhK;����cV���t�+��Nz�+������ҏ�` ���1�n�>��d��X�ٌ���$&3��Lcz�3�f곘��2��,`�{[d�X_�Roz�\�
V��լa-�X�6�����J��6��#��N����a/����6��a�p�c�'9�����g9�y.p�K\�
W��unp�[��w��'��2��<q��|�s^�W)���ڼ����G>�ٿ�%R|M)�����'����?PK�z`  �  PK  ў,J               147.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=ÇW�&��:�b{{�����kW�R�~+n��;e�K���+_�k=]�R��[Y��Ȧ���F'��y��dm��Y�_,�J��X�@Ol��e���B�G:^nO}k�J���}�y�n�>d�j�ҜyE�|��1��_2�|���Z�ǌ5I"煑q�������I�{�n���N�e��{�������y)���Zl
�0�Kcâ.\�yݵ�I�a��Zֿw?S�'���i����үc��̸�*Q�R%y���ɧ�m�9���m�5-ߺw�b�<f�t�x���焵�[�u���=B|�D��'Ei,ڢ����~�us���jƬ���Ur;�m=zr�ɳݺE�4K��'�'X�T����ti~R�n��`Z��2FW� |�=��a�oKzBV*���*�Yj�y��G瞬2fظ87�u��uqB7��\�N��m�%�5�P��&<�o�[=�ÃL���rs��r�mg�2�$���X��<?r���0{��nK��?�)ָ��X�D�\��"����M4Sn�~�.r��_׽eݳ�o&sV�����Y�{�QbG�޼t���}��������T�P?�쵗צ����հnA�勿�S�Fl[^������/O.-����EW�c"���p^������)�7��~�i��i�|�B���8�S?^�`����ua����ŵB�\�&Z�,rUd.p�_��6�����sv��˙_3닭^4���<��'�|�~m�͓�s���~�_tU$�g�t�|�YNu�ic�'����l�ؚ=��v��S�qJ���r���Y׎�Dn*OV��i����/��_{}xqq����������X�����Lsl�B�K�){g|y9�1sZ:�N�������|�[��;��*�T�u���o�dNB-o���U]d�	te%TJɾ����5���Cq�CS���W��9��K�j_���k�)rS�O���]]��yl�}.-h��y���7�2uq�$Z�v^�~�z^�S��r��`��sԼ������u�ƣy}��$���k��l��	`(8�t���	 PK'Y1��  �  PK  ў,J               147.vec���Q�wv���]��]���lA��Vl�V�[�V�V,�?�S����=?�7"���S@!E�(Gy*P1eQɮ�^��T�:5�I-j�\Ա��ף>hH1�hL��4+�fzsZВV��mig�>+�zG:љ.t�����3�E/�7%��/��� ��Av��!e��HF1�f��8�3��Lb2Sҟ�j7M��f2���a.��|��B��%,e�Y�JV��5�e���FJ��f���ml��vȝ�b7{��>�s �8(q�#��9���o���9�Y�q�\����U�q��������]y��<p��G<���e<w�B�L�J����|���x�>��]�)��_�7���J�PK�eV�f  �  PK  ў,J               148.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=ÇW�&��:�b[{�{���u�A[�̄-[��_���a�^��l���/���kΛls��r�����2u%��2Pg�.�lz��͟7u���zn�v��Tjf��D��o�w�3�=����{�҃����Ϲ���U$t!�K�&�t<�y�9Qy����v2�]��]�ʢ��7�Eڪ4'���B����h��"N�)7���#�cd��짛>������e�>���]�Ѝ���ß�Ԟ�Ǟ����ͣ�����pi,j���e�O�&N3�Za��d����M6����QO�d%i\�9ؿ0�^1�fu�D����X�@׀�.�Lx0�����l�vM<q�=����1)?�߷?�[��ٓW*�s��gk-�x�l�c����\t9 t0>���%˯��ܫ��%���z4%1%��Mx���ǫ8mT<����YO��̝~�٤���iv]�]E�`Ƌ]��������Ž��H�~Ƀ���lu�v��
O74��dx�F�ʓi�s�~to	tem%�����mݾ�J��&ᬄ��'��˯-�S�1-�]�%i�܍ ��v�(wR��+7n��4)�����;��ĺ��X�Zp����e��?\}��I6%p�������z�gȼî���I�s�Z�}>^�f�+���&Ը�*?I�覃_��c[�>4�������5g�Um�x�Sbk�-�a�r��Wo��&m��g�ܻs����a�*������������
���x��㸔?�����P=�Ţ�T|!#���~��yj��sF�4\�u�����W&���8�@%,�(���gq��#�+zN�P�~>�!Ù����qW|Y���c�>�Gw���q���F�Y̢.	BQ}��w��S\��o�e|����o춾ا���{���\�<�?��T~yW����^���"ѽ�F���b�����v�^�J������}q�Oe�nV�;�e�-^,��7����s�e�2���7� C/'Bo�d\mT���e�fݗ'N���M�n��.��v�W�Y�㮸����nq>�r��Z`.q������ PK���  �  PK  ў,J               148.vec�e�a�=�z���n�vv7��-�b+�b+؂qU�[�P��������2ÎȲ���(�y�R��THYT���W�
U�FujP�Z)����u�G}АF4�I�h�E3�9-hI+Zӆ��K)�g��w���BW�ѝ�=�|��M�ҏ�`��d7X�P�1��d�m�ȱ�c<��$&3%��T�i�tf0�Y�fs�g3_.`!�X�����`%�X�ֲ������Mlf[��vv�씻�������`�7���(�8�	Nr*+���g9�y.p�K\�
W��unp�[��w��'K��W�P>�1O�*����U��k���
�N����g��%R|u#��w~�_�N�PK�>��d  �  PK  ў,J               149.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=ÇW�&��:�b>j�i}��v�9�N카f�^�w����9���j�J������yLS�D(jڋE]	"����9نm��߽%?���r�*�g9U8/{��{hٝ����������*���B3��4V�h,�b��_�ڞUpq�R�2/U����_������3M�KZ�MԈ=��=�~��#�|��-bN_X1CgהK�&���x.PT���@��d��Yo�jY�d8ab�J.�/���-}=��D�g��5��"80���'��6Y��D-x��4�]��~�u��x��[��o��l����A/�B�'D�[��k�Ƣ|�jo�1�Rc��������8�Z�{�q���_��-�T�����h�u]j����&��wlv	fXԥ�3����T��g�U�"��ߦ�d0�޾r��c:�4�v������t��9�����&�D*�d&}�K��r�����W������=�R�?2/{���Is租�R�U�������kM7r?J���hb��H #����P���!�==�;x�x��_�e/�=㫳��J�U�j/�_='��u����:��_^.c�搟a�0�j�f��Ʃ3
/�t���cmۺ38��8"7#���pٕ�.���-�'1g�ɥ�EKui,3���ǂt�)�u`E#�rK�3���F���t;rkR�4�i�Ӎ�.:|�z���]֫�bd^��>�Φ�O�ڽ��_Ze6��8wɦcI��nܯ�"�oo��b�&+ۃ��,����zʻ��WﶖKӜ�?er�ѵ�	J���D|�/��6�ih�zYt6���:v���#���z#�c�c�^<PQa���h�|�u�v>_����xR;8�߬��'�1sf��o��	E��ڡ`_q�����y�g�|�F_%Pj�9��q�_sP/�*��H(�+׮���0ǻP��A���	B��g�>W�>��K'�䈻��>e�U+����a����Sn<h<`��z��&u��u�ˊ�[�yo_[cg�pC���� �//}�f̜f9;�͓��{k��o?�'��S��S�ړ������X��7PK�X��  �  PK  ў,J               149.vec��Q�wv�l]�c��ε���l�[�[�l�Vl�B�Q߮�G��s�f�Y��
)G��T�"�R���U�Fu��AMjQ;�NQW�G}АF4�	MSD�� ��Ŵ�%�hM��.�����A�H':Ӆ�t�;=R>zf����}�G0�A�c��}(%c8#�(Fی�c�x&0�ILfJ*��v����`&����2�f�\�B��%,e�Y�JV��5�e��� 7���la+����s���n���}�� ��8$s���8'8ɩ�,N�3����E�䒼��r�����[�6w����=y�<��y�S���s^�W�v��ȷ�+��{���|�3_l�F�o)�w�����7R�PKJ�wUg  �  PK  ў,J               150.i��eT����P:��A�a���k@:��K�K@:��$�F��������n|������:���y���</<�T� (�  ʿx^�^```b�����|��	.6691>	5����������������U����W@@ �"*)�'��/���MP^�|���C��K�GGE�����n �i�7 
= �H��� �;':��?��
DC��|��_B DE���������щ�xe0��-0��H���^0�����L�1�[����z����������]@PHXDTL�����.DO����������������磯_hXxDdTtLRrJjZz�����¢�Ҳ�ں��Ʀ���}������ٹ��ť�ͭ��;�{���W�n����� D���?r��BEC�a����?	�h�t�D2ژn��|�/Hd�jz^2�뜑Z�Ob�b�`:����߁����/��͵���{< ! 8{#��	G�ˆD-Q圇�C��B���ο��*y���CA��sKG�mbӁ�ܯ��>����|�Be�m���V{���R�4r̥���
���nw�~.{�^Yx����kL_	z��BN�['��|:̳ڡ�%�  ��:6����sG�Y��-%(G���V>�#���������A�A�_\w����s��v��r�V�2вz4QK]��u��(�eGK\����	C01w���\#B����0���=��F���_M�1��?�AO5��Ċ��Y�"O�����~���@���k�M��u�Z�;��W�gJ���y
Y �ȵE��槆q�g Bs�!-���ǃ�f�Y�.~�m'�1U��3��(e��Őw���QF�O*��}+��;o����t�������f4�s�����u�~�3�h���Z��,�"��\.��&YE��;����8E���8�*��������[١���ё� eg��z$�|&3�ܬ�����X�7?A�B����ԉ3O�7����d�ª��Z=��+��t��m��2*_�E���3 �Q�j�Q)Ss��"̓��W5i"S_2�������J�_VP%ln%4�j\Ǐ�abw5
����䢴�&k�~�	�BF����P��~H�~��!O��g�9H�K��Q�M����U��9�-i����=]�6��e�~\�s�7�R*��*^��Bw�r#�%��ޘ�����<�f��lRyA�ĉd�'9:��M�7����`���v�� �̽��|�Z>i��,���V+�DZP
�Qy��F����p���|�x��+���B�2�]QU��O��Dw�卉©��XQ�BN;�[+��5S7f���80I9��P=�l��$'�N��#���3v�Z���O���W��ѐQLq2^��^>r�[s��&M���6M�r+��1Q�jxЃ`$�n�aq���`�~�ŕ�P����M�.�]҅m����+BqĜ��Cc��LDf�'mZ�"�Z��=���~��;+�����h!��ȊE��jB���S5��&!SҮ&1k����_�������H�GƊn�)xY{L�����)j.>-��� ���qR_v��Le�F��;�����<�l������I�ɓ!�
��B���E?$L���@���3�?yJ|�����^]k�����Ͽ	^�xCʶ�ѽs[��I��Y��obrfV�d�,����6bi!��ݘj#��g��0r�;w_�$�V7N�'�r]���J��35��U��s����e�HpIS�_�"vV���M�m_�<v�V��N��Cm�$��T�����75;Ղ��Vu������'�j�;}ңc�S��]p�3 <��Rx/��Cy�c	\�̺Fn�\�}�s�
-]B'�E9�k��INi0�ި�BXA'�H�n�Y��܈pt<��]c8�Vl.MX�����ah������J�_W�[�QK8p���y 싟~�MU^4 ���o�[s:���˴	�8'��R��o(n���_�6j����Jy:��|,�H��>�A��Y�#�M�����㷍��Ug���-�xcV�DW%�-aK������_�y���u�C�+�5K0ȍuD[މ�X����H��|b:&6�3������ �.��t�E��}4�d�x����.W�nP��BI����ʝ*�i��+��ZϳZL~�\��jn��2��CB
$|��\f�Ye[Jo$5ef�N��0�ǐ�����M��˟�#K%����WD�c�L�-�Y]�9R�рE�c�y�H�P�[���R_�
Sp<��Ƙ�}܇ӛ�?j��zk���#��{U(6����TO)�o�(���GHC7Ua�'zK����?�@_pTwv�ƕz�e�-p��y�������b<������[�>����*���%�g_�bb\Zȯl�'��ai���#�/�����{���4�����4\.{`�"ϤL����VW�I��Q����|� �٥���Y6G9�m@�C ;�tN�3V*��� �����5JQ���9�^����G�G�܌Zݰ�O(e�hf�l����5��[���V�LS��� ~_ɘ��u�1Kޕ����C[�����Ay��픹�0!�%)`?S5KG�ud���6w�n�K&�!� �Y4O�G�%��9��h}}W݌�[{��In3C�޼f�M�R���qԃ�sD*�~/
��bF��7�`��|�ە>�s�$��жb�|P�}��kTN�� $��4�T����7�c�lVz%eF`G������	�YKM��@��ܾ�P�rO;<62�����3����˥�ɴ� �%S��E�R,�qᚧ��w�$�`O��3��0��9ҁ�Q�F��������]b�o�v��X"1_���1B�*��t�A;�� �85�?j�2 &���/�cv��b�u�S��j��������N���	���Ie�%������7V�����q�څ����ixќ�ٓx*.����s�4��Y��*kLt�I����zhk���49u]��Re�Z�xF)F&������JE�%|��ZKrսZ6�(�#3�#�G�oJV�>��h[�ߙ�)y1�����;OD5v_�:��e���h�������7"��ѓA���zt$Xv��5}����M.{�2�
�T��,H���F��a��m|(��Fe��{M&�OM	���W��_�+4�d$�k���y�4Q�����D���z�A+�Q��OP�$�u������bl�'�s��Xr��!X�k7mIm�䜇�m2������*ܺ���Mq\~q;Y34���8��2�G�$㉁�Y3+���FJ�t��#���'���\��H�����~��Q�)�o:�'i
C���v��hg�a����G\��)��yrt��]��;��oҝf1.�ؓZ_*�<l3L�^?��&Tfg�ǥ�;/`������z=�zo�h�$~Wd�6B֊tDJb�h84UY=G���
��]#π�ʨ,���:�삩aE9���T��
��b�S��bD�"���o�ݵ�޻��>%=@n@�%F�j�Q���-"1��ԁj�P`�����s�(�@S6�r��@�Z.��k�<����M��
uLB�4ʩ��� ��j3h�=%(��p��������e<�k�]n����XAg�_}p�%��M_HY|�i��#��K�7`���b���*>�s�̙s�)����r������l:6����2_]kyS�.<P!s�p��x��O���&��O�h0]�ʝ �s� ���GG���V�f��h���-P*�0��rsl��/P��V9�X4��~t֯ş�G�\�B����<��n����U�xD����X�����ث�%0�I���<є.MIP��?9n���c����)�����ECѕ�I��@�����JN��?�(n�$K��R�e��6a8-k��� ����g �U����)Ҵ�kH�sT��G��GW����%)_�z�]����0lo��Q�K�Y�p��-�����VD40#�d%�n�ծ�x�㹺�߹m�[�Of&�(H <}��86P1)�G���a�6�^(,t��Y�����?P�zwP�D�L��l��X��Dq`/f���Q�T��6�Z��GӁ�)�a���SS�=nF<V<*�xm��"��{.;�ԉؖ�6��x�:m�����d_L���>^���8,X'�U�}_�a��ȯ����۳{3�:8j�ä�DPw��t�����I��-��j5'*��8��r�|I��ɍN�
�ߔ�Z��2J7��e�r���6m@�;��ۂ��ǧ�Z��=GTU�/-I�hv�2U�:���C=B����ళH���ɵ�m�����ܩ���y��fYG� t[[q1"e��yl�e�X+��
nR�ܿ!jN�WK��e�'�������:���e2PY�}�/H����<�!d���k�2:k��y�������Zz�Lƭt�r�CH��w�y9KF����DLaC�-c��'�%ESg3���S��O�D���v���I�o����aMx0�
��&%^���+�c��ptw�ϟ)��	����/!�+�o��di�=���_�Zy@>�U��+M�&�+yܷ0������U8�$�cu]�!S��qr�[y�G�@Ș���5��68Lkm�e�y���fn�[a{�����!M����E���G��
�q-�
��'�	�Z"JB���ǏW�-�_�+�2	Rx��Zm���P����<764o�T�_aEr%>F®�\WnԨ]�	�r�/�BG�&����MЇIs�EǼ��G/�K�!��Tl���~�ȇ��D5d��-tZF�Nbc3c�$3�ȶ��(Z�M�%U���1�M�q��"����9E�׋�U�
�Ο�
�s�Fi�W^'�2Jߤ���q��:�,l~֧W��lu��?���U$�T�K�˾z�#���ǭ9W��d�36J�|��2Љ��45���O�{e�6�/.���]AG�L�H#|Ų���K�"�g��O�귽�ͷ�bo�a޼��
���:����T�O]�o������W�l0O�z������sB~3�Ff���ky�����y�\���ȸ�R�`5���x@7.�;��0+j3٠�ު��Z��`�q��p��5�A��4oG��B���7���?Y8U	�F��`�EФ��v#�FQ�Y��'�P�� �9`p�M�=��{�MBL���k������D��ux�,hI���nũ>��Nm�:A��;�B6=�5a�d0���?���ɢ4׹�1�kA���zjN[�L�
����b���F��$y���%���"��؇���1��5>"�i�mlc�@c�.���Y�6h�Ae,{T�j��d�;/�¥�c,1,׌֕PM�*���hoSN�̊�������R�]�0��9����v�6�T����R?�-[�,�z���'�2q�V)��<J[S�_7\n<F�"YCr�{ѓ��M��q���衵pޘ�䱻,1kNz�&�(ڴc-�#]�I�-��!�p��������j��'X�T�,���R�����N=��of�Ԓ|�q�ۯ���q�*>�/���z}���Vʍ����f"�-���zo3�vt�a���y����@���X��~�y�M���3�y%��I��8P��^1��3)n�p5��6'.cŧ�4�%�[�6
z���f�w���cu_ȫ�xCm��םN�>�Q�abf��ͅ�̜f4y�`A�_����/W�'��ᘽy#�>ߢT�)�n��h��kK�L��m#�s��$ݖRZ8�S�Vx�!?x9ˎ�����}0Q6�@�,"?r���i�*��D���wӚF�3:d��88���F���j=����I�5���J��]:��w��J������JR͛�Y�F�"���5�T v]�;���҇ZW�j��C�9����� U8����`ڡ��x����[�ݒ����gi��q���NA�l\�r� ���E|�q#� �wy�p�X<s(����c{���Z����Q�H���Z���:^�(ď֠��K��0��pB����Y^7��$'��0�s-�zuq��%�̀�&C����Ҡ!�R�k��\�5#*�d�Տ��"	�I�uE�؄��� +v�!HB��C�y��n�ԃV� Ȉ͸J���W�P��p5Fe[�����=���,Z"U�־��^�ݎ����5� ���k�U9-���|�PE�v0��)�J���Gj��%�S��x�W�1��`h����X�P�*�:�z���*<��7��0�VmSPw��W�肄|�9�G��=�Pى���,�#Z�	���4|``&��Q���$c�Q���I~��l��9Z�?�6f�����DeZ������y7r�L���� a��n�d��i�Wjv���|,�V�eCq�Q���T&�&��	�]@�?� ���L��~�7���f�rnB��G��
� `�`���r�	Vɼ��l�$��Q�$4��_jǓ#�b3ꈐ��d�������h!�.R�A��K���g@��!���#��'"�?���ܖ�ܣ�l���%%%d�>�m� ��P���+P�[w����:���� ��W�a�M��]L��а���`4�5C�8���O)��љ�n�r��{t����V0�C�>[�-���I�#\R]e!��k�G�s�лp��խ��J��a���U�jZM���㱷��`@�l� ��.�*,��Ѕ��ƗI����(�m�5�K���,
F����"!K��!Q�8��!l���{�$BQPU����C��նh�4���b�5S� �R���,����e�����Ԅ�\�˒G����X�[OpӐ�LA1�U%R������|���\����S�-�$�t�%K����ȼk��aE��@*%+�;�st�:���O�������o^�ƍ�� ��M�`V��ל�R��?�|�p[���I/E؆��F7��QN9C��H���>����t�-�����W�TÞ�����Z�'W��[�ݗ���@[�CF�+yfP�Q�ҤF�4�hB&��VG�95�S-eW������N���x�+����ce����Z��բ���T2�8������E�6�g���TQkB�'���+��)�'�5��(�z��(���aJb���r��fP��[�|��)����/�tT6�r�����S�"!8&��K痏K'��Hj���>!j�!��E���^r�Z���qE�&wMei�����	kЊ��	� r6�7�����i�oj��)�A���q��~���=�{f��L2��r���M�8�3��2U�U������k��i��W+[i�1�A���FGtor�7Mӌ熤e���C���;�t%��_���C��D'�l��&��x���lO����;xn�c��TD��X1�[���WJ����P��u�wq��枫�zٶ
:���:ݩ{�C0BE�45+�oO� ���u> _�Gv1,y-����%��oL�8B΢L
Rd�p+�ָ�&�`����i ���4���&O���w���QB���u7�>O�ׅM��"�������}���s���4kk���ZB"ɯ�}в�Z�j���{2�R�b�-�u�u!*�SuÖ�f3�ws�?�Q ���_�}�}���8��f-�S�8r�D���e�%�[�N9W�f�D �u�&/@E~,�V�N�=R�~�Xe����'0�cg���u?���xd�s���]@g��
����ݬ{@^B�e�S<����
��xUX�H[�s�%������M�@>���"H/2�W�N|Y�����O�?#���>�v���Zʘ��ˁ���B��&������l�p�t*��&w�#ph�)>SXH���K�MW�m3^,�/}xi�����<:^�g���U��M��e$�o�-4�� -���"sSD���Ofg[�+δ��5�d���m��]2�`�]2JJWc��W�2�8�9��D�|Nܑ��![q�鯽_�s��r��0\R�B/���xu�yy+qy�N�����2+����hOo��r���c���m�J� £"$�z�?�c�$��&F�Oտ���TT\O��az��I���j���a��U�0�o?	�
7'���[߬TzLIi����t!���x���u���=��H�x :���fyB����4��:J2MZbv�����r�(v�mf:b>��m���ҏ��mJ2Ű�4mOB��S���k��R�!���3P�j�o�*��̄"�ܔ ����PKxb��5!  �!  PK  ў,J               151.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=ÇW�&��:�b�a�Y�Ħ�M��m��7{�$�����AVo�-�գ��b���%���_��'���,�Yԥu�KcQ>l57��G��'J�`f��gu�}�����g��^vz��ϻ�Ƿ����\�����:��²�4��>5���'���`��^�o�g�<�C�>U3����r�l��'�jtsgXui�ta���e��ܚ�S�7%��L㤛����~�u쾝5��꒝���+�+��?�c&_j֌7�{�C]��40��|�����Y:5����)2�c�e/ͳ�]߹Fa�{ӳ4T���5���{~���C�:��"�!��4�`�%�FϹc�;'(������iכ�ٿ������������J���pŢ��B�z�L�(4oM�H��Bf/�(��ٺ2�G�O���)��w��Z埿������=)马�V��5�_=���}Tv����W]���1�_u6����	�����ҏ�Kʢ�L8:����*����
��n��f���o�G��%�Y\ �'���p�9�k��پ��rr׻-+��9�M�z�g�n��/��m����y��ooO[*T�j{3H�U$X_X�(���ky�Z��D�2g�_��)���+�#�lf'ܟM�-,|��#5����;Sx�4�<��j=Soi��NuѻΦs��nr�%x0��y���F��\f۪{�U���p��I�W�k����N����E�(�i�oz�G�d�{Y��Xy�*�s���}��#G��4�y
�?�Iz"��7�kR��?�Y�9Ru}qE����&Lϋr*2p<���u\�Ŝbλb+uqr��[�z�Ni�0y�.i-"`��������Zs��/��yn���u�����M�*ٙ���f�>�H�F_�D��*@?�h,�b@ƍ�F�3�P�d�{8K}��?u�շ�
��L�|�������+u\V-Z��j/��k�nuG߈�X�$�U$����� PK{2Uщ  �  PK  ў,J               151.vec�e��A��=�cwwww뵻[�[�[�l�Vl�V,�u��K��������,��'G)��S�2��\ʢ�]�"��L�R��԰��E��kS��ԣ>hH��خ�ޔf4�-iEkڤ�h�E;�=�H':Ӆ�tK��壇ޓ^��}�G��@�A�`��P�1��L�e7Z�X�1�	Ld��ߘb7U��tf0�Y�fsm���,`!�X�����`%�X�ֲ.��z���lb3[��6���;��n���}��w<(q�#��9�ɬ$N�Ӝ�,�8�.r��\)dqU^�:7��-ns�P����y�=��R>�'<�y&�󂗼����w�����G>�/6_#ŷ����O~�?)�PK��ٙh  �  PK  ў,J               152.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=ÇW�&��:�b�a�Y�>��=� x~���7O�J�`�1.�.z�U�����;��<y>���N�+W\��κ�8*��A����S7�┐��r���ꋾ���ȽL��e8�]8l?���g�ϟ�f�<��U$  �U�f����I�E�t?yp>��G�#O��;���[s*����iɓ<ҞY'����늶���s6��?+⾮����u�N�/�"��*��Hh|a7ճ�!�2�En�R��0�E]80��;c}8�j�l�xw���?�;&Ⱦ���~̬7�f�b�d��j[���ϲ;'<[�w`�Ƭ.�U�LD2Y?wٕ=7b�*n�8V��㺈g��Fӻ?6iL�̵�VDa����I��U.{��F�����H(�Ƣ.|�e�{���c<g�����9���:�S�Uo}T�g�z����ω�ߔvF/�f1�jy���W�$`����XԀ[��gX;a#Ͻ���}b;~�WO~�����y�>���o�>����i�{�Q�Ibo����r񭏾w��.�=���XV������kK��4L_^R�Yqk�ݣ�1��L���'#ZP��m�m~Խ*u�Z�`R�$̾�J��o�g�v��w��y�Q�z�w�k���O���>��$�T������r;MV�;�5�Ţ�T|A|�k�6��o
��������mv�Qf9�}��N��Y�W�i֍��/�m�-:-_˩�]����k{���*O*�4���F��kO��7q�gx�|��Ԭ�c�u/��	te��Kg혥+ev�9g���ׯc���	�ߑ��b3�fF>����{����ЎR��/��9�Ô���e�T"�M-Lq/U0�� v�����-���U����p������An�#�s��=<|��!Q��A(V�oU��V�W�7���3GR��}.�4I�6��R��y��z�
�h��YqP�r�ʼ��o�Q��h?W�,WP���J�+k+Z���^�x}a�sXނ��%
'5�0w�����N�s�{��;w}K�<��)��$3Tq��.̮tU��d��7PK���#�  �  PK  ў,J               152.vec�U˕A��=�cwwww�gw7؂-�b+�b+؂�؊�X�?�(�a��ž��Ȳ�r�)E�Ҕ�,�R��*��De�P�jT��]�,��^�:ԥ�i@C���Y>��MiFsZВV��M�m�B���Ӂ�t�3]�J�T��v=����7}�K?�3����S��2��`d��(����2��L`"���~S��Ә�f2���a.�����,a)�X�
V��լam��ur=��&6���l�>��v����a/��os@��9�Q�q���8)Oq�3����E.q���y�k\�7���b1�Ȼ��_�@>L�x$���|�s^�W������|�#��l�%R|M)�����'����?PK��Gc  �  PK  ў,J               153.p�{4�i���3��Ǝ�Ȩ��ĸD����F�La�l�2��"R�P�R��z�-Z�Bl��[�2R����v�ٳ���?�}����9��|��}$������v�v �  (=�d��$�B"�h4J��bde1x%ey��:�KMuA�d����V�@ ��]��J���6�(�F�T�R�F�1�5,V��MЦ�cIjE�H��: D�*���(�~�@G QhYiC� �P
��`�j����J�� ��H� �/����Nűk�d�ɎD˨~��W�[�O6XM�hbJ33�fC�nkǰ߳w��~g�^�>�|��s��	�6,����b����ˉIW�S�7nf���),*.)-�Wܭohlj�������ao_���gχ�GF�^���_ψg�̽}7��P���KQ����0�	YjP���7 ��0�A�:�3(�V^zAZ��qJœ�%�J�>ӛ^B�H���"���`p ((}<�"`L�Ȃ88����`,�S�� �|ΌwlX�Q��ޢx��0οX�6QR�X��4Ε �����Ѡ�<zK�-��%�A�Cc����Cj�w����8ݻ4��:�Z�ı�5Yzi	W���k�"αI��J���^A�H���Cs���-<��?�Ys�+^��.9���G���A/U��j�#ƻ���;Ϙ�(%��!����ۼ]E�J*{��f�k��|m!g6ҽ��uk�α�D�a$@���u-�5%
��?��hD�6*���x��db�-� ��q�SI�.����y���c��i�L����>c���h �����{�h�.�4�˽�rv���r�O�B�X<"D�GX�.�[������s ����9}�w�,��ɤ�ɏh�p��dUN��A�R�(��c�ֽ���o�-/��s+�7M���	��=��#��G#��������_ԫ��>�-��iV#������OE��	�71�\�Ӊ�QFM~�q�}QrϮ15^� ��hf:���F���M�4	p`�u����@6���k��cҁ��
M��y��Mc�TL��7y���;�M��ɉZ�%�4�4��8=�&Ģڤk�>$>w(���D{h�p��W�[��䘦y�$5�Po�q���Ȳ�l:���n1Ý�nZoF�p�8�U�I:X�rC�MÒ�Ω�&�e>��F��*�U1����Z]D�z;�L�WV�W^-fx
�|a�ӻ�$@�m*'����=�-�G�*���r�c^��ϫ����;=�8p#����g�׌\^tluT��&���TʫS6Z�u��%@4�ҏ�l<V��R]�N2[��+&>w=n�ӫp���E[@5����Z�FT,�zf��ھ�{Id�0�h�ic_�bB��UW��%[ލ��ۥs�Z"��X���?�1�%��fX��,k�[�blQ�q6�|yf��%����kWml��$��N�����};�'���%(�ru8X��|�L+C%���;yiQ�\kv��W�m�!2?�R��WPKJ��  �  PK  ў,J               153.vec�e�Tq���;vwwwvw؂-�*�b+��-�+���X�j���.~��꜉Ȳ���(Gy�S��TJYT���J5�S��Ԣ6u��f���i@Cј&4�Y�h�EwKZњ6����
�1�G'wg�Еnt�=�e�ۮ��/��� 2������F2�ьal��8���	Ld���T�1=��v3ݳ���2��,`!�X�����`%�X�ֲ��l`c��M��b�P�V���6;u���^������a�p�c�'9����z����<��%.s����kz���������B!��}������}�e<�y��x�^�*�㵾�-�x�>��6_"�ה�~�?����PKS�0c  �  PK  ў,J               154.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=ÇW�&��:���[VC�}�4n�������dx�>����Y���?��R���'E��r��_�:�/S�H`�G��1��U��g2�s+e��]���2�s�ZZ���<�5׳�h��T��'d�?���7\����=Kw���	!S����m�}�Uخ�^%|a��[k�4l�t��c��`i?��������Zi���j؊'�d�6�Zw����	L��8sc��ؾ���öGU|wN�jSt����Ճ'��~]9�8��j������{d�+:��z,f����lmY���I����ȜW���f��5]t]��*���'���,�B��@�r��?�-S��K�5�mȷ��M�>o�� o�����i��pi,j����xW�
�x,�{����_�z�pf�W����^�]ֺI���(���ơ��j'�ei,Z��ǡ`��>���`O�f�������v���N�n�n�����s�k��I{Ʈ��-��=u��������Ϳ������g�p����1�'E<�u_�`>߲������D��_k���,nQ���H�+>��c�w�ʜ]=*���j/�_='��n��W?�^�X`��t�Ϝ��)Y�}67��"��-�͜"w{z�*�������:���|��׫�����xkޣyb�KrN��|{e��y��e�r۵��4��ƽ'W]���40���U_��W�g���m�>�t�y�Ӿz����l��rۯM����"3��v&_'���ݒ�3��>s���_׋-g]����w�L	>ƃ�NIs�����.,=����_�o^6���]��O��,��8qNf����\��m�[�%��8Z�P���ZW5�t�.6B�]n��v���0�E�<X�7��W���z�a\�z�ٶ�O�Vv몐�������؞'���
d
[)�bQ��a�r撍�[3�u��q�j���6��h�L�G{��Wߴ�=g���JNK�7�/�l[fMj�x����_Ş�f�Z��3��FW��6L�����'�����GNg\�U|~Y��ƍ������d�K��%m[zJc�X>a� PK��p-�  �  PK  ў,J               154.vec���A��ww��kw���b�ݝ`�؊�؊�`�b+�b��QW��p�3Y�O�"��S��T�b*�Jv��*T�%T�5�����E���R��4�!�hL��4+�fz)�iAKZњ6�M�h�壽ށ�t�3]�J7�������7}�K?�3��6��`�P�P�1��t�Qv��1�e��D&19��)vS�iLg3��l�0�y�gY�b���e,g+Y�jְ6��:��ld���V�y��r;��n���}�9 r���(�8Ή�o���8��r��~�y�K\.��"�r����&��](�y�{��S.��<�y*����U��k�����=��'>�|�_��w~�_�N�PK/��na  �  PK  ў,J               155.i��uT����niI)iXj	Y`Q�	��n�\RB`�\�X:$EI��X�$%���s�����}�;gΙ3w�=�9s�3s�g�W �:�� `=4��@@��O��GH@@@DDHLJCFJBB�@EMN���򔙑���S��������G�9�����7PNJDVPTL�?A����HIH����Eؘ�D���@I�� ���b`Sb�Pb�wX������������O@HDL򰠞���������������p)�؄�u��]hD��s	9�j~����5w&"�{L�������9�����PZ��
XUM��o }c��faie��������듷OHh����Ȩ�Ĥ�Դ���¢bTIi���Ʀ���]�=�����'&��gf��W����[�;��'�g��.���Å������|������%���P��	�S)���P���(����"���Kk�:FL�)����?h�M���E����7�<����p( �&J[� �>A5XF!��I �_�6�(��+x���T.X'�6����S���%Q�NAM��r�:��6�&ͫ�ġ�9.���u��=�z�X\�����+���ߔ6�|���(����$#8a��}\�e)P���wB�/��Y�X�W�������i���af!�~2��ŧg�@���k�����NYho�l�A�
���&`�1��MA���0�����f�Ev��bL�"�=�g��lR��0SINW2v%�1�,U
��2��-� }��b��mf�oed��kbM�9N3�z�����~|=|��ax�-�Dl����˓�Sb�u:i��9j7�[T�*�~IB~j�j6U1��/�2���.zO�$��L�(�yz�kr������ŏ��@��|,����6<<)�z��K�6���<Y�l�����<�x&'�m<����b�y���D+��Im|��ѫSP����g��.�,7^wuE������! �QF�f:��^~�O ��(_1]+�u�w�vbnA����7����0�i�s����k�+��
�ҭ{�`r�K�	bY�	�,�@6���$�x�1��-h�� �s�bۖ��9_W���e	c��TA�᥍R[�;?x�`ou��<f�5]�ɻf����	5p-�� \L?o5=�yA�qJ7���g�Yq�/쵣��k�'���'�kD'-�s�p�*��늘����i_?|ėP����v� ����U�Ů[��X������m�{@�]�l���!��!RL���_$��z߭�� �Elp�;&P�Y�~pFgM_h���ӿ�$�Y����#���ci��)%�B=}�]�������ǣ���fT���M�!��1�v]��+�y��Bʅ�E��b��gt��E>�좑o��(O+U+iy���em�$Ⴗ���Yj	)�
]3�vv�ye?���q?^��M�Ҡ�j�����6�)�����A�=_�QIDVV�œI��?�Ń�J�776������X
!F�O�(�;z�� �U�9G*�(�{�!�,Ҧt?��WQO-�K�؜E���hVf�W�8{��6.�9Z_6�'*^C��Uj^��(Ia���&:X{��Q��;o���M�G���O�B�w{��7'|�M�|vϪ��/���_ed��;����璱��;��]8�Tˑ�\�O��쇰tch[�"���̴�X��+��|��;>�-���}e���׋ފ�g)4oc��W&Q�;i�N�4���l��U0K�����*n{����u��!�:*�9Cr�8��Ǝ�!GC���.������2^V��@�'nw��R�h�]�d�&�K,��U�kTG�?/��Q/��E`��KB~Kh������s��.㱁u��KR��b�����������C�'��x�����h'?i��hW�r���4E���4�|�K氣G���8F��v�5���(h��awh�~�I���=��Xp��8��x�HE��2@�>�j�`���C�7�}NxnG-_a$�P-j�͘6���ss�-�9~��"uВ�L���	�Y+������D�f1�{x��(���Q����\؎��$�R�o�i���NmJ5��m��S�$-�υ�9p� �Vm�M�˴�߲֣3�Qk̵���p����j��|�jz��V~a�k1�Z�ٔ����o��=ϝ!T}�����W6� ���� �TQ{�^�_٩������@���������S2=�W�M����� �$L�u�Xׁ,�,Ŭj�-�A�XCB�u!`��E��2�l"bE]e�I�%x�:�2�K�Xo,��p!�Z�B��ZW��-,��(�E��ǂ���D�&���q��F�lј��J�.m�C ��tᘥ�d�Ȓ9(�u��a��s֏�~��v���棆r�%w9������A�?`@?���)����#��{�Qs�h�����D]����d��|�F�i���e0+R#��D>7|q\�w�)e�7-�	�'Y�Z����QR��!I7�Z�Y�9*��x9�?q����Fb�mc�Y�p�컄l�r?9�_�-W�{'����'*���?2��p�D����ʬ��j� �-���o�3��!�sm���	��X�n��w`�$2���A���*ݷ=�T��/���f�R���@�yXE����6s��5��0SF'R�&K�^dO ��d���(���Na<��	_������	�*���ހ}9�x����c�_<R�w�-B�bX�Qv�Y��x
T㫭A|d�ж/�<ͱ�x)�`�foV����U��ѡqW�����E��̶f���s���wn_Y�MW��?\�#�w��9[R�ƕ3�QЎF1��P_'�ȍi[�u�����։4��P�1�Y��틅�å��q8�?CV�DA�b}pF�L3���\nj��|��kNU­�>0���H}����Qu�s�A��\M��û�Xˋ�P_���ip��xg�~,�/\� �yK>'$]F��.��4�Œ�)��S�}������2"���ӝ��OtBd~�pJ2T�]^E�q#�2���A�Ֆ0z2��}�J|7Z�/�5z|�јz���e�n��~4@5`����v�FUO��s�{���w��-��Ə��9ܠ��Θ�>:!g� ��0��WdL>��.���,����"#Ƌ{�Td�m�B�y���Y�R=���K5wpa����pE���>_l��w��=�n	�W��$�Y���|�S��y�ն��/oj>�WucC�g)4�!wH����4�]�;���Mg��]�kB��"����:Br�.O���Lr'���!Ґc�V?C+_=�.�<{��}%�%��~j�ĸ�|�A&�:rR�Ļ�6�K\��^n1�I?^��k�a-o�I�{[D�����s8��o�ZJ\�	��6�2�J�l�({�Ѓ���� �㾆��7��_�(Ou�T��t_DK�X?nʅ�NO'ɶ�}��-Gĺ
���)A�$}�A�:DB�o�i:9r����=y�3��?��U;�M׶@�'�f)�v��o�Aݸ�0�[]Y��<���	)T��vM��s=ݖP��&�7a��m1��^����`;F���Q2����� :P�qp�1 �j�K�B��Y&V�1�H���y��� 񜴳�SI��I��p|�KM�����*(��= /���ͧw��n��-
�G,	��kM*1#����t����X�?.�m\c���+4�8�b�M��jV�&|��RAW ���H���S8$��&k&��j\���二o��̆�:6{P��`��i�J���_��o���t�24�
Ȣs���\C��4e[�-�r�"0�'e�6�j�+�}�����p�0��R����G�/Zy�k\���:C��+��8;^���]� ����6L�Ă�:�cf�3ڞ��+s4w�K�=���Pg�P�P����������v�4C#sؔpf�/gdG!��<{k<[�3^09��W+����i�Mf"�1Ӆ+aoV���뇹�J�X��5�����FJ��Z�|��V��������/� t��Q<i�J�+�b��r�@��z��_�dC���3}��$�[�	a��&�!���4*��(J����2��l�����îƏ��X�3UDz�?q���L,�Fg����3��3���e6(�����x-��b�K�9w�RXQ���j����h
e��;�˭��S�_O��,�E���\[첬g�+��l=��yUS�DG�5�m��>)��D�惒��F$�c��r'���
�	�|̋��z�Q���>�(''=�7�XA�n!o��k
"eg��/VΆl�hm�͕���rp_\B�R�uu[D��5��x��?�hMȶl�6IѴC�+�Ody͟���`=SOT��/	o3�4���e���Hk��/fNe�s�j�Y9��O+#�}��fr?%���-uxT��-�r�7Z��,vC��)����6"-Iz�����f�F�J�p� qx�A�I= ��^i���(������<�D��Q�D����}�4��0Ա��Lg�e����j����%*$*Q��8q�, 0�����GT>����?�'�U�x�//�#B��((��8ѺAgO7-I��c�����6��,�q�U@%4:����{Y?Z����̅eg �t�<��,%��%x����Ek��4>�E���	)��"-hR7�N�	F�=��h*�&����rK��,��t�I�= 1�Y�D+���@lvC���Z�|�tx��>/sc����R�l�N�Λh�_�v��Q�7�4�r������ӏ_F�ժ�֪�
k�Ym����Y��qF;ӂ�p�["V���OK���˦�ϭͰ^E*�YY�Y�CV������x�\�&�$q)�P����*�*�6N=����0� ���O�0��!��T���ag��>Y��N�d�����d��[�C*�̈�G�}[K�si@�Ż%-*��8�$"���iwvJO�ۖ��4lF'q�����������c��Mԟ��~ar�kJG�����zS0�y�.��$̠����	��/d�:/d���ûDs��|�#t��K�������HR�x��02�I�`Zrwgٺ=5p4��bn�u�n,q<4�n���`e��Ҁ�O�K�S�ݯK�׍�f'���_[`
&�B$�?�\�d���k��{p�V+�)s'	��2|(P��O\E�V��q��H�Cv���k���vGQ�{¼�s
E�.����7�m����D/ݒGƫ��8��Ǖ��u�z�M^C���m'(����k�p��3~Pz�4C��m�|�l3EՑpH/T�W?AZ��]�L+B���Ŧ���r32#�����i��l�Z�IqTZ/�A�����x?NNɥ"Y�v ����e`)ⵋ����ql�OZ��	e����c/���zA��z�YD��u�4V���.��0���~#%Y�U��:U��	�+e-�4�:`�B���� :���`�qz �m
T�z4v^���ʫ�?FR��Z>�gp��n�7�b�d@��'����sN7*M[qr/z��8�UrB(��D/
B�Du��&`�h!�4���R��z�R��(��A+��^-|������*>�kک�Ǖ���3������C喴V��>n�n|m�1'��6D�z�m��1�T؈r�cUf�v&�;dk�QsL��ٖ�v1���e��U�]�N��Mƾ�:������c_��B��r1mƬˢ�_�8s{WȎ^GA7R�˞��s�!˚K��i� )���ҹ  �d޳��ۯDZM�@N�`m��6�n�v��o�� �#�M�3�#Wխd�J�ѭ�D����(Ү���\��PV��ަ���F��������W��ד���"4�<j����5g9Z�"�Yu/�Y� �I�t[���5 �+ד�G�)�ה����4s�/�'�|3;&��{����,"ɽ�y^�~gS�c#a����7�T��&[����x9�Z���{բ:�>gw����6l�$fl{,���'n�*R�L����:2�䃧�)ɭ_<���DT�g�տ_\�6��y٧�<d10/��#p��e�0�k��v+�[�L�B�;be|[͉��N 2P�}�!_}��G�)5�@p\~�^rW�<�(�0,��	������v��[j��:<�x��"&1Ɠ��ySS�L^�Cͤ7�J�s��%i�I0��$�R�W�U�1)̖b��u�����񎠕�?�v�XqAk)���,�����
Sw�_��P�Y�K�z^�JЌQY��K��ܲ�������n��j����y�Q�������|ņ�8K�jVE�gZmz�5�=	��͔���J_��٠p�%�[i�v|=�~]Uu������8~��ϧ;[hW���Q�����LQ;=��;ɓ���G��A��+��0�ݨ>ԫ�����K��]-�����#n�c�.?d���J�0�&�N��'��(DM�ګH'���{�ʔ�I�����r>7~9�N���1�0X)�W���9\_�?�ʤd����&gTj_"*��n���#���e�r2%.ȕhX \�H��'�Uk��.��f�2��0Y\�����Ɵ
c�ˍ���69�i�q�̪�.h�GD2A���HL���R�DTS��g��hQ����Ru/Kd���S����6]���3��^ϗ�_����T0y�"%�*�隦�sUg��y��5���
�q�5�_��&�N�D���4:cː�]#3�k�Sۋn::	�z#哱+k&��x7ѵ{|A���*��qos&+"c��Ū�o��e�=��=#B@���y[�e����|�п������Mj�c犦x�N&	r�p����˯�����x}kZ�ά�΍=�,%�:'�J����l��e�.��{�6�_��=p�/���Ϫ�ݎ���vN�e�igw����$%�{e��+meno���q͠�yQ<<��n_��uk>�σ��U
��{�W�C���!���}2�z�dg!_*��*�HX/���9��?�?��+&{:���]T�RY��n�oaZ������7KpR9ҩ�V�Yi)�/��_{���H���?�cO�Gq^׷��1���_,aVТH�\�,�	���Z�6��5B�?�M�e��C���?�S366:��8��ɵ��c�t�D�R��x��x?[D�8Y0��-n|�s�b��5p�'�~p��|�7�1�^�YI�Ä��������vuZ �D|l~�N�]���r�]w��@-��`�tF��.�e�͓�&P`�����R�8P���s{b�ݼLMo��&�nK .J��y�'�dug�}A��ټ��Ⱥ͹��2�2Tl��h"ɹw>a�����p�y��mË����uP���g�n��q#��.3ܳ��e���T�,K�N��pc�,ĸ�������/�у���
/���q�1K�,�+n�M5Z������=x�c9�2�����֚mΞ�����,E�J�ߡ����7[��UA�����]6�~�g�����Zf��A�~����4�v9(��c��JS��	G@���U��6YkF�f���5r�1!�����
���(�l�t�OQ���
�Q]5��'�)����'AW P!�����{ (��7q4�8Jd��3�r��7ˤ>m�	�Į�,�������iN"���yS�x�_���%hd]�&NY[4N�h�8���j2����Ci)S_�r�gM곿�p�]Լ�D�[�C�{��O6���!u ����f�7^�j�>ϕKs���	i ��bjb7�ɝ#} �G�ώ�b��#_�\;���?.�6N�]���p����~~mU�mT��������>>H����̈́��ωJz��m�a���0QN���2A��5�bE���>�D���FAt�x�mf�\`(��1�9B��= FB�5�(?{�a,�I���aFxUsd�ܷa�*0{�JP�OJcG<	�</#G�8��НsߊF%7y��Em�/Jl��́�T��=��K@&��zΦ��>P`���FΩ�痘��f�AZx�+�t"�̓�/��w��QG���%e�>�Q�3Q�E?Ħ�/1�gͩ'����ɐ
���p���rR�%�GuD�Y¼���?�*��*�t3���~���Q{�9C�w�\�n	�.�Q�3��WN�`���.r{�H	��̹Y��S�5���Z�IB�̝m���\ɟ���<���B	d�r���99����ce��!��K}L�=`JG�\e�MDm�������C^�5|��T0&j��-�쿳�f�6����AO'�ǝ����_ ��2V�-�Ƭ��!��lSu���ʷe�;+�o#���FJ��=V��n�T!u�_�w4��z�|ot��a�7�c�_�JZwh��s�PK�/�B!  �!  PK  ў,J               156.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=ÇW�&��:�,�ܚ���j��j�(-�{[=�Ns��y^t���陌�E׽���|�xK�	���]�E�]�f���k�S��&:b޿^f�wYf'����7��;�㉱���,{zF�!�U<���v��m����1	��?n/KS�2���.�QY��ΰ���^�#�ߺ��~zf����o���S���~��VT:*��*���G��=�m��H��}bם��u{���Q�LO>��Y���|���'�ο����wmV�s��=8�t�����6��E�z�wk�콮������ۿ5M*Xz�n����ui;�\��1���rd����-���v�K�QY��L{�G������� �*��F���/+y�{�Y��\>��,�����V�.�����XW+�/�-��ӻ���ĉ�q3T����m�}�������t���@���N�>�U�։q�B��I[�ݑ��f[�����E�5'�l��j�gz����)�-�Z��辉\ԥ���������:��k��'���<uSOo�g��&�|���wV�T�=�NR�m��q�����?�r?(=ДH}�/�b�A�o>���41XX�����1��2��3��;�m;W�hj�]�'�(��|�(n���:���^�j��=�ַ�Nso����j��+�K;��z�����_�hA��O�'��hû�S;*�����N8�tr�܉e+�-�<���Eg���G
=�'�Y}U.x�����g���$�w���}��Ks�H�+.�Q'[�C�+��o#B׮�����r�΍O���_��1��d�m������W�,��>���>?>�����+��JS�7�%7E��z4�������Ew�Q{�@���~D��.c1��-<y^�>ƨ����V.�K���~f���Ʀ�
��?����*/�X�afP#�,N���L\7^Ir��wg�����_�[����M\�?w�+�����"�i�Uŕ_O�\o�?-��q���U��"��ͯj��qg��m��q�+K�]e�5�����ʍ&��}[hr��S�˓�~��[��Ə���W].�z�ݩ?�س�gF�F*0�, �c$�d�y�,�H��?CɃ����Uۃ)9M<��0�����"ɖ�E�'�~� ����t`��b��o PK��#  	  PK  ў,J               156.vec�e�UQ��x�����c�bww�c�-�����`��b+�XX�?�l9<g��}"�J�y��sT&O�R��)5�,���Ԣ6u�K=�� E4�"�iBS�ќ���]�,m����=�H':�%�k��nzw��AOzћ>�MY���` ���2��6#�HF1�1�e㙐RL���Of
S��tf0�Y�"f����2�	ΗX�"������`%�X�ֲ��l`#���[�V����d���n��}�����9bsT�8'8�)Ns����<��%.s��\�z�"nțܢ����.�
��/�G<�I��S���6/�K^�����o�k��{>P�G>�/|��)����7���?PK/;?b  �  PK  ў,J               157.p�YTSW����H��X�
e4��TB
�e	"�	�Z �����h�
�"D!������0��aP�ʬTEъAd0.۾8�}������k�_�(۔� M��N  Pu e'�@#�($�B�0�����bqd�<Qg��:�(=#3c=�9�
��d�<s&��klm3���1��`08,N[]]��O�g�c)� -4hd@� �!-P)tUs"��>�Ap�ƨaU�5A08�@��*_U�Z���"��ʀGd��
��<�6��هQ���6y�l�1̈́����j���Ŏ,�%�K]V��\���^�ݰ1pS��Нa��#"���| 6.�� 1��D�ɔ�̬��sr��]*�\\"���U_�����߸y����-�m��=�{�<�{��phxD1�f���4@���(����Cp�4���G�#	��(?�F��pL\xch���rWm��{��4�{�����������A�*<H�^��2D����3Ŏ\z$�V�ٱ}�sB�a��QR�"?+ltK�q��>����ЋY��5�Kv�z��`=y�~J�#q�-S ��G��8�Q3��`#��
�	�X[rq�Ǥ�78����3�ܗ=Q���#����Fo=s�%c�S+^��7��2�D�0J��6:�� չ'@�x�2��]i�&3�H�D6�������j�T'��ty­;я�h�j)�X�7h��a���GPs�_�:��+��D�P��
2�F$�~��~m�{D9<�u�J@Ƚٽ�����`��''�Y$�>��~�(o��ԜJ/a줸���6pDB]����b�ST���lo?�)Ņح�Hl}��5��"�`���3�:��ԥ���V����x�����������7�^��)���KX2,�H��W+6��>t?Q@���R��iei"'������RӤ����$�乕�E��^�7�����)���a�-̦x��b6�Kͥ=Β��R���!��#���o_NA�tih.r��ZF�m<"D��hKj[���ؖy?�� H���=/���r�锎��n�g�Dq�����Y���9�6Ѯ�Q�jӐDв?δ��]�,ny" uį
�=Aw�ߒ�!O3��.O����Rj��ۢw �\���b�*s�Y��6m&���⌟�PHP�	�M/-��{SG�����|r��p�3Y�)���ޒ���rm�lc�������D\���ӷ�)SXq�Aj��
eA�*���+-?y&�2z�?Ahl�:}ɿ���!_}׸8U��XM�X�9�ۻ�ͧ����^�>�,S���μߛJø�{���KM���>�h/\���������oY
��6Q���W�|r� �U�ã�A��-�3�����z��k��1�k���-�{���T=3�N���[KE��jO���X�w��6G������������xJ��K����{{DU�����K��,��M.�M�лb��Q��Υ��k£K��m��'�׻W}$t�Y����<�.ۘ�&��1O�=oDw**N�	�>xRБ7�
^v��r����l�PK�n��-  	  PK  ў,J               157.vec��VA�s]?];�^um���\��l�[�[�l�Vlŵ�P�;>ry����\��ȪD���.�*9�Q�Bj�\�̲��צu�G}А��(�h�7�)�hN�iI+s��[���-�hO:҉�)�Y.��]�FwzГ^��Oʢ��~z0�AfCff��HF1�2�0�q�2ƛ��Od���T�1�����L}���\�1�,d�Y�R����d�Y�Zֱ�l��&��-le���Nv9��r{��~p�Cv.G�Q�q����9�Y�q�\����U���q]��&�ܞ��w�g��|�CY,���x*������W��oݵw���|�#���;_�W3�"���2~ȟ��7���?PK\3��f  �  PK  ў,J               158.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=Ç[�&��:�,�p{��]�ٶ�y��S~g�[��	Vq��rr�^ʶ]:-�g�v^�_��O�z"���q�+mٯ\�QT�wbX��*�@W:bƋ�
�0�����p��\O���w\Sh�����:���9����E����m���_̵7�3Ǌ��|Nm��_��Y�����oS�yN<f��Ȧ�B���w����2�l�W�h�.�Ƣ�\�pa��e�4J�:���/�x2�8a�����k�w\�M��V=�{����m���Q�T~�������ݽk7��-.z��u�I�^��۾�
�Y��� kF��&OW���V<�&����␿:�J_^��8Ƨ�hk٬����R�^q�K�L�gzL(*������"�������b�V+�jy؇�gx}������ű��:v�BUrt2n��y�'{j���7W��,K~��k!>ǂl��U}Ϯ�˷g����~��[t�=�P����+?*�v���?����j�/�e���PW���H�c��H #���K�o~��������ʶ3���ױ��>��J�)�|�.u��_�)Yo^�����SN殓�b6�k-g�u�����;��]-e��+��h��+�fKW?��4Y�.d�)�E3ui,`y�K)�w�1��]����A��mB����q.,4�h�!,v:yY��0��9>�~߲�٫m�����QB��J���ϧ�9��/��v3�}�Ub������,Y1�sB��-ǯ�Ox�=��si����4�t�$�]n6�5{��şx�+�5�թ����~����|��-�h��-���֍!M�f~�l���Cn����k�L�ظq6cjÂ���?�S3�}�n��7��>%쑏T���N׷:�`�����^���"/8���7��wK��|г�������t�E,��c�w�W?�.U��S��v��m֍�/��y���1��%Y,1��'�D̿3�1��.u�璿��
��L��R�����Y	�з���>y,�T�����"`1����V7]Q���~�����WW{<V���?��.���\��0]h]ヾ�&�.��s��Y��K�	3I�Nc�\����Q����"Ջ�00�6,�����E�'m�B�����@u1��	 PKq���  �  PK  ў,J               158.vec�e�VQ����kww�ح��]��`�آ���`��cb+֨X�?�U�K�����Ȳ�
(����L��\T���נ&��M�R��)�A�PoDc�Дf4�-�Ze��ZoC[�ўt��S>�d��w�����'��M��E_�~z0�AfCf3\�`$���2���oL���Ob2S��4�3���6�n�>���c>X�"S�����`%�X�ֲ��l`#�YQl����V����d��[��c?8ȡ�O�G8�1�s����4g8�9�s��\�2W����5y���zn��ܡ�����y�C��x,����|�^������w��|��m�D��Y�o�;?��/~��PKy�kUa  �  PK  ў,J               159.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=Ç[�&��:�,�{R�b��=��n囩����ѩڻ<-TĎ3���?�3��b���JqW����3S�T�[�>���]/�F�H����H #1���),�r�9I���V�d2�Xw?j�]Sw���N�WW^�,��P���k��y�5?����	�	��K�8/w���s�&s����}��`���3�<�ᩛz��
� ���/�t<3�4V1,�����7]���ib��\��yu�M��&�fﺞ��X��z���j��7(]	!�ȵm���j�c��F��?����*������oVR��_��?�{�.���6��G1�E]	"���p��殦\ק�W�Ny,�tuG`���c{¶���u��y�ߝ�
�9�W�N4��[ԥ�ť������w��?C׻@�ԗ7��������O����4�{I	�{J����8:g�?;�8��.	tem%�:���mi������~�q�ﾏ��{>���~�P�W�a��W���~/��;Iy�H�g�<C�ě�ghM�b�}�ݴ#�l~��/�}�I�aɳIᖕ����F�gز�e�w~���2��4��j��E���j���?l��S�=��Qу:э��\}n�	�g���X�%v��e�)�yb�<+V���R�v�>&|�=�������<�;�e�������&��Lg���?�����K}䞮�X4_�bk�Q�󱃋?��f��Va�4�ڼ���z=�&m�?01r����{��ݪ�H�)Ͳ>x^v�̉�α�)�{�ދr��iw��/����?��cL���"x0㍊��o6+ET��k<{�O����������T#S.���{G�\!T�ٹ��/���Z����E,�2uqJG���U��<���ќ�:��M���������yKo�{�Ҟp�Uc��'�M��snr�uQn�{�?0X"���-���e�z�^�x�������%�*V����=�ܹxc���ˑFg�'�͔v-�u��P�������e�.J�0�Ţ�TBŪ��� PK��  �  PK  ў,J               159.vec�e�UQ��ܙkwwwwa�ݝ`��؊��
�`�b+�b돺�Gk�^��e���QD1y�P�r�O��`WQ�De�P�jT�5SD��8j�u�K=�Ӏ�4��]�,M�f4�-iEk��6�]���z:҉�t�+��r�î�ދ���/��� ���B	C�pF02��(����2��L`"���ߦ�Mէ1��d���\�1�,d�Y�Ҭ(���`%�X�ֲ�f���F6��-le۳��!w����a/�������9�Q�q����9�Y�q�� /r�˅B\�W��u�7�Mnq��y�{����#��'�T>�9/x�+��|�[��|��m�D��Y�o�;?��/~�'�PK�kd  �  PK  ў,J               160.i��e\���X�$��n��ZP:�ZZ\J��\���P:�������|n��/�g^�|��w���s?u�x������ ��~��������@��`
"�G`2r
Z#-==� '+==�3n>A!QQQ�$TBXF@DT�?�`��������际���@��%�b� �I���X�� ��9q��� �ð��8�x |�Gj���@l ..�ì��< ���YH�\�-�řB8 &�U�F�3|�&b�H@H����������GTL�������J�*�j�z�pC#cK�w�6���n��?y}	������������_PXT��������������ή�ޑѱ�ɩ��յ��ͭ��ӳ��W���� �����H��qp�8��paa{�g).���6�39�p >�BL���UD���e���Mt���?h�M���E����7� �z� a�Ħv���^	K�% �g_���Ĺ�{)i�K��jW�#hZs�Qc�?XT��u�`�%P�Ǘ<�֋Q��n.�)�mP�W��r0`	1�
�`ᠺ.�ε�06K�	-t�MF�k�Kj�����tt��cE�'b9�wQ'����"Y�1��!���J��u��3��Z��*��]�۹�<���W��տ^ ް�l��|i�=+|6L�
�t9�ߜ����/���JZ��OC�^Õ�}�ۛ8]��j�슫����������GZ��UT����h6o�e~���|�"�
��n ��(�`��#�0�5h2�.*d��IXi~�t�Yu���m��I&v�v�c�M>+����N
��DN���ԍ��9�%�vi���N_�kiٮ4��y��$�eL4�}�j+`-�]B1fV�cj�4�;�F$YI�;XG|%������ʛ�iz*M���4���_0�]���׉d䛺��tA�'2�ʒ��k%�h9�s����I�}�h��ǪF{�$ �\��i�t���WAN�Vy�!l����Z�(ЌE�B_yHAd�$��&�R��k��ƒ�Ǩ����a�F ��T���p�:|t��&Lev3���H��s�!p���yG �#���^���?���񃝹hl��Kb��8��ɪ�w"\��ҍ� �zʞ_�̥������L9Rß��N2Q�B2������[vZ�i����Hg��)+,�Ź�Xޟ�>�V ��`h8���o)t4��3�����\"�(��A��V�����#HVaAM(?eo�Y�����I�$Nd����N�����Y��%T��7^6���cR��ņ%Z���W���M��Md@eo�?1/K<ۇ����;{��灺w�S�J���&n�s��m
H�-���z�6-��@��L+%��*H�"�Q
����D�u�S��d0x9񛚃�8a�I�"���W���|�;R��ˑ+Ƀ�ԉ<�&��V	�L�I�{�Tϸ�Q��I!i�_0��D��-w���[���˼My�t�,�X�P���9^[.狓]����ԁ��os��=����.��_uG�^��^�Ϗ�h��J�P)���Y���k]�Ϣ�M_�S�Jٽ������;�x��8���T�<4���ZZ�N�B�٬/?}ի��D���r����&uj �&�cU�p��3�b���c��%�ti�ݿ�ucye �����',�q�.���nOO��F�;;�xE-YO��f�C�4dns���ζºG�0;|ʺ<�pH�%k��K�(��uF��B:#*�� ����0lEGXX-��CT�w��F���xjl���6��b���\�<�zD[Z8�n���t�	<��"�r=J�s���#�$�(0r�S�ʲ��Vw^~��J��߫����
m�8BIN��9^��ƭ��)�=��Ů-e�|��E�<b��ka�8Yg��8��X�lڸ�L=5Ӂ&Q�n����I�d���L)7h�倞�7��t57<-����'��J�g����������+��rrk}k+��k�t� ~�H�-��[E�(џ����G��2���.B�ոx�/�V���g����X�n��@�b}�8�1y�M��7JQS�11@k�����g�5���6pJ�zi�`����+닋�>�n��~G��G��Ƹ��_[���+�}:���,���a��>'��n���%�����x��J=��:����5�#�+=�O0t�D���]���6�Y"$��q�d��y��'���GX��Z�Y���r+�jr��kGo���7�#/��2���Y��T��c�ǒ}X���	!5��8d$�&��u��]����]���d�C^	͑G����O� �V����y����pd�cE֭�裺 e�+�l��@��gО���d�yci�A-��]�W��o9��Z�h[ͧ�'�Q�Ԇ��t�ܬ��+7��K����]#g(G��t���{�d���o�]�>]B]@������V��?�f��b�U����3����|��Bm�n����qU���}gk���>���.�0{���p����ST���=`򓉨�j�&?k�����_M����f����]2������-8�ѵ�����d��	X�&�r'��	*/���nw~��~�X[�oپ3�o[
ցVi���K�d�,[%��փn�k��[M�u�nھ �{`� eg��a���ő� �+=�g
��(����;�m�/��H2�6O]cE�^��9\���94@��sx��ѥ����=aׯa�a�Z�yq7�U¸qÖ,�?D���ѐyS�.��X���z��E)"6ƹ0��-_x,���&$�U��+�hVԸLr�F�)ڠh�'�Wj� ������:� 㶈?��<G4�Gޮ\��w��=L@��b��i�́*K�2ӷ���P�Jף����sb��&�&��.I�� �Q",��� ����k�l!�r�J)�[�2�Li�0�y�!{_�o���@4O���Ӟ뮳�=^֧k�&j۩k7Lv�1:0g����7��%�H�z+��l��ƚ�t����>���ޮd�Y1(��V�Ć��#����5�:�#G���Y��$�#�l'4��(�7�
i<1��+�-��0Vh���v�ִ�+�	iL����N�x������Ad�ܬR�&���9�=�\�i�ߕ���!��C;�U5*����-.�B���˲����lF;2�f<v,�A�~gLQ�8*iC��b�дm����x���s�L��u��)Ma��d�����ׁ(�͟3��~b��p*���	��>x���6�]\S�[qF>�@��V�{���	��g�%�D�H+�G�@~��v���h��b%�S4�o�FMX����&i} �-2�w�~;yL�ì<*C���c3���� ��������7������Χ̃�X�k�;a��Hr�y�̠�3̓�`����Ɔ(�Mi�`v8�]MF;���ֆF*�xEԿ��</����@��4����^Y%��R&9a,O�Վ9���!l��w�vF���k��0�	v.(a�h|䊂ޖ�M����ќt_c�vKcxy�,1��3���8���z ˆ�L�ô��?��,�fk?���<�s��çڛ�p�a�'�u�%o�#m;&b����v�= �~GX��
�&��XeC?��{C.���ߑX
7v>�Z<��O���[�`��4}�2�7HA(m�pG�6�;M�0�ˊ�|���`� t�7���%�N���5nnTo3G��Ă(>�`	o�GG��UC+�NXr����U�g�5�_��S匢}�ҡ[���^$��IE/
Q39G.��Ǒ����Eh8O��Gq��I����B�Q���/D�,�y�ֵ���V���q���U>iڼ���=�h4�T~��j]�`�ve��*FNO� 1W6b{����h�Ӓ��O������oڐ��|���9eJ�&��ղ/������Y������)
gӵ$~f�>Ѝ��2ރ��8���k���ѳ�g��ٳ�?�(�K+�&��&4�ʙ;B>��(9�����)�5��!�pw�i	�A�l/ݨ�R��4�����z:�w�L��-ڹ�<�DI�,�ه�H�@�o\��S�H�ئM$ �������Φ2a����@�Q7w
mt�B%���3ؖ^�i�G ��u~�w��=��.x��7QE��W�ݙ�
9�j�?�l�I��%��'�eG�8�ר��E��J�ߜ:����'��*�[�9	^�(J5�RAo)��V�Z��\ PϘ?4E�J���~��<����^�q�]*�bQ�_*@�.�T����>�;�w�@wg�Ѫ�/(����9�������k��.紻mW���/x=bkU���E-b��џ0*���O�㤖�8K*�=�A���Ѕ�=4j��"	�(6Ui��qw���q�<�ZT�\�5�m�S�BN�%{Ag��랯U
ʅ�Y���2��{��B��`�O����~��Q�\!����I������&������)`�OώA�';�6vL�B�X"���O�w%�5a�U�e�ۿ8�[Bw�|s|�(�k����BuE�&�R�v�f�:�^��S�2�Z�#t�`��ߖ��Ԏ'���~�0�u���o(��an��TheD�tl"��U�ו��"���gNU���y��U�4���Q�l<:�p���zdX�3a���J�йA�jD�ո�e��`7j����ŀ�|�_�)3�ڗJ�Q�']��{C	�4[�HAC���i��9*���y�}���4$O�S��3���~�M\�u`PB��;-QR��I~KH��HX���KAǗ��mK����Q>����5���Au0ƺZ�W�
=y��� {Փ��FBҚ�*j��H��z���mf�#f���
������7��.k�t���jK�#G\:�0�O���{�ރ��5�q��%�(��O��5��S�Dƾ��h��j���j#^�����/	ÞE��\"�/�1�,�"������ut��S$�:���Yۻ�Z�On��$Sؿ<��^Q�h��wٵ.�i��{@y�Iǆ�C@]:嫹�HC@WH����|��̬q�e�=�����	��G�<�y�f�Q���2�vɶ���t���?���L�`�af�;�;��B����PF��=�}��W��������V�`�]��-�q6�W{^u�Ŕ�F�� ,9��ޅ� O%A^�A�n%��t���Ğ��v�s�6t,��RW>v�(y%QJ#�3<���m=�趸ݴ���v ^"�V-�[oy*��e�axه.Bժ�I`�;�IR}w��Ifs�M�e���PHR�����5�:u�^ϏeT|/ë�����ϋu[ހ���<�vtII�	����Sle��{�ju���֤_a�=�����ʗJ�}��*f�Тc�2Bcҩ������/џ[��6{wQ�s�\e|^�w�]U�����obA>^ex��>/���U-��RDg���&"��$Ew��?=�}۽�ꬨ���ϩ�ۛ�߰w�ׅ�U"�e3��5�W\����y�UZ@xZ� ��`��U�Xɫ[>��ZEZ�F2�m�ڻ��X��t#/�cqQ���Jz� J��_vڕ�HА�q�[W{���;֊c�<��S�����Z�(����ݺ����,	���W]>�}����C��F�}�S8�PPTgv�C��3�K&�x�������_H���C�7�ԎF��xU'1�2*X��u�9,�<&s��}�7�e��2��*M����L*�k��lGO7�T�����c���g�������W=�"�M�eѯ��?���٬[A����*��/RSR���֟��r(y�}l=\���Xs�"�Y�6��F����{r�d;���R�q��^��dx�N��G�"�S�z�(�zt��Q�ֽ�c��Ҩ���9��ȑ	'��/O�K����Se^4U���N�����XP oj��O5�wL׌���ލ��6���Ҁg-Q�Ȅ�+|�z�/�6>Z�r�n���?A͒���mCi���/�b;��O���\����}�5�_����Y�|1>��(:E���<eK�g�Iq=�DI|<n�o��J�BA�|F�z�j���ζT� �K8�Y�GQ��zM��E��G?|�US�Խ��p�@Xl͵�Yn�Ƃ�@��H�Pct��+`)=h,�0����0�uϒ�Nʹ����)uFܸ��6�~�� �ӈ����R��A2x:�ҕ���s��=�'��f7M��(qd��'r��<v�O
���鍗������W��d���/�}Ƃ;��h�NX�}|o5�?!W��E��s��4��Eq�o�U����޾���q�M�.�'�����wB��7�y��RMtpYD@����TS��%���O,�c�A�>���Q �餃���i�j�L�[{��-:��4˥m%��V�A�t�.�E����m�Nv<���'�g�p4��b-���0+�|�D9)ن!�V�אo<��{�p�ZWD!BnP�c٬��<��9T�9��%Y�֡l(�:��A�cY��чp�=�������]4�<�hӸQ��l��]'b���1�����s�����\��|I��@0_v������T��zвJT֕$�[�ǹٷ?�K�!��(nr=�a/Ȗ�Z�{]��2_��n"1�p���X�i (*�A��/G���q�����1vIW®�5痸�h��bq�R���R�HԲ�'���AY��D���
�S�|����>�������>���ة9�X�{���	���v�2��R$(͗g�����`Oꕛ�²�'����.X��{�9{JAϐ)���̂})+��z��x�UfN%r�F��"X�Wσ�+; X��Z��+��`�Cɣ4���}���C�>�Z[֥�I�W�u��^�����9�t���{��c��G���qQ� �4Ֆp3�sc��pL$����5�g��_J����N�b7�?�8�j��r���/��J���9��M-uV�k�nٍ�2u��9�	��M~͖:y�3�y�ɸv�ǩ��'7Ύ��	+]���O�����Gkg=�6��./A%B��X�^؏�Fx�βl�*\�Cf8�����CE�*�e�g�
�}d��Q�-K����Q�g��}(���R�KG����|ӳ�j��%��i��cF�y!��d��C��Ԑ�hmE
0��C~�4�����
����7\����DR�u�|)��+s�"L*�V�E׷��i�ȣ%��s�۷�ꈤBv��i	�Ʉ]��̻��g�[���e���1�Ra)(O�D�F�ݗeJ��;t	�-H\4y�u��*U�,���SF�&jo�~��ȌC?�7m���^�M�N�(�r���̤��۳=�7,�c|��H'q@���^�Y��T��_��mOb��^N���Ø�V�E�ae����w�kj����]������A�t�@��5�"O<c��nyg�7���gb�
�9�s�
gR�!>�U GWfr��<}D��>;���݌�9��P��WǙ�k^�L����aZt`����찝���l�@i49oa�x��{'��t]������P�w%��톞�T�>G��/}�ύ�V0�:�n�W��Qǐ�&G�f���]��6�p����b������=`��_��SGb�`����<���ݖI:s��#DuȠ�&��A���lū�`�+����dZ:�i��Y
8vj~��&7����;��Co�_!٠�OO>��6�v2O+��w�H�Hb���<��b{^�d�$ϱ��sg-�̚B--����|ԡ���8���&�˕[@�-G�EK:�z����C��qs��A����+/�\��Ͷ�>h\����3�m���GR9N$�3���/�}�1�F����c�D6^Ţ���֮��Td�8c�X���B�rr��E�Wj*�X(��S��o3<nv��]�3�O�K�74L��;�0&;(��
>2ks���9U�H�c�y,ƴ�~��f��r-����^l�;5�'��;v_�e�x>����!��R��b�ٜ<�㍛X�v�0x���'��oX�R#Z�����/��{��TҗB�Ei���%J�h��q��Pɜ�������L���+;90��d�A�B�����E4�C�Z0����M��ǠЭ-�$v�
�=�4B�_�D죂xX\4	�d3�ȠD��+���C���Ui�2R�l�����|Y7��/r��Q����9�8�&�}�̳��G��ݟ�#y�Vƀs!��l�zT��ugl����PK�#�   �!  PK  ў,J               161.p�{4�y��w޹��fB�CF�Ҙ)�\2�R�HYr��ĸD���2e�v
M%Bn�=dR�!
#��RrWd͎�^��������;߿��<����瑴J~[s�8  P� I;�	@#�($�B�0������K�$e�*IYEEMc����UE��N[Gw��$k�36��c2拀��).Z�Ƞ�P�X�* �M�LT`x@��� ��] �#�(4F+M(Y�@��!�FK� � P֘"�p�Q�ADF��Kh�Ya��]㈆��(FFa�����r-��
&k�:}�����K+���;v:��������w�_pHh������b��8+HH<w>)9%5Mx9�J�՜�kEŷJJ��+n߫ݯ}�����/[Z�ĝ]�=�}�oG��'&�>~�����C˅�r��p���a���pe�`�E�-QgD��fg/Vc�zv#��Ff���<���;������K� P:<#b����5�?X��J���WˀU��y��M>XC��O���Q�{Vq�1v���BpJ�
܈\6�_8�w:��yU�rr������vVsP�.���U���,�Ip`|$<DN�Nvk��h6϶aw$|�v�r��>�U}9h�W={=���z�(..�P=4��A+�q�|s��ȏr�m`���l�:���3�V�u�G��[�_wɿԗ�̄��R�;�ж���0��Z�z%�˖���	#���a�mr��Jf��5��	���EN���eeǁAq�Wm��ú������t�N)�O�\{�Mܶ�Q�]�v��rʃo�<���Ӄ/��tѵX
�C�m�*���:(^fT|d�;ѳlM��2��eQY�M�k��D�K��^gW�+F�O��Y\A��W��ϖ&�m���J�n�
h�����Zfy.Y�inh5Y=W��ec�`���(�_8�讣k42�DӣF���m&��z,=>�e#b���$�8o��W$H'�G@���ݓ����1��xBj��>��_V77��^���c��	�C>�Y���]ڱG�C�5��1�mos�e\�:۶�G�)w� �1�3�8��;�3|'���l�g��"�/0 d�)�����S�q���Q���=���>��,�'��+��ec
�m5�l9��@���] ��;�=���upH�����QRc|�.���'>��`�F�*a��hB�5��w`;x�yMW�f���%�l��]7�����n{�����k�í�๱�v5�|�e_AD7G-��1#�X�E�U�=�܋:��}�[T/jxȌ}m4�0�A�Ȫ?�B�	c�����ƀqO?��N��!��UH�(�$_�@f�k���.��Y�cz���n����޺�Z��,�y�̸s�=�:;�����yM���B�"j��w�QG���	��%�L�*Q5s�{T^�w*6��b�����¾��:��F��:���CWU%�u��'Wz<�7���M9�)m:��[�,i�PK�0���  �  PK  ў,J               161.vec�e�Q�w������]�n�l�[�[�l�Vl�Vl�Q�����a-�����,��O�<e(P�r��B�G�,��^�*T�թAMj���Y>��u�G}АF4�IJ�Ԯ�ޜ���iC[ڥb��
�A�H':Ӆ�t�;=R.z���{Ӈ���?� ��rC)a��HF��1�n�>�q�g��d��L�Ә�f2���a.�����,ai��er9+X�*V�������ld���V���?�!w����a/��ρ�4�C�G9�qNp�S�.fqF����E.q�X�+�*׸�nr����Ȼ����@>L�x$�O�3�󂗼�y-��w����g�/��k�������'��͟��PK��f  �  PK  ў,J               162.p�y<�y��9C��`���ϑ2&G%"4���jȑ^S!ef��)Q�q4�r5�E%���t��fG�=������}���_���~��s|%��g���� a  J v�
�F!e�h4##���c���J��Z$m-"�L3�#S�t�D�\�h�	�� �YZY�W�2�s��+�%���"���Mr�ɀ6@�0ǁ��$�	~5�Wap�����I� ��a8�@H�l�@��J�U(eW?4���'� �c[~Kŭm�f����UU#�k,�Ճ�K��-,�٭�wp\�tr߰q�����m�ۃ�w�D펎����t0������S�Ϥ�M���^�˿t������j����v}ÝƦ���u<����{�?0�b����ɩ��3��@ �fʅ�r�8=��b�p$������R��d��/���蘺���G�ɪ�}��о��=��E�;�\� J����h7�KE�]m�R*��Bo��a�\ ��ޒ��OX����I�B(�7�T�{5�����A�Dp�|���!�ȕ�󙀳A����
d������ �O;��;�b��~�Asb���"W{���o im��$ך8��:|F�q�Ӭ�w��X�7�Ž�s�LD��*x��F��K�3�J��J��8b��[d�����.m�B�S�IǶ��	�a=�ۼ��(��J��#uդ<�_8��5h����蚁��Z2N,�De\��ܲ"�]'�y]5v���I���K�{
MI��柿�{'�]�q������將1ͣ9r�(�T~4�bʲ�qC�nՌ�M�P!��Y;{���-�i��O�']�M�Y<k������P�;��:N��Gt�ԺV�
���d�A2��Ҟ5�����mJY��xW��<w��+.����&�a�k9�G�ɤ����s�͋��946J���Ӹ�;JR�W6n��� �̧e�	��B��P��k,_&V�>6��Y�}�S�A;D����|�S��S�E)G��E(��2t���M_͗�?�x�|b~F��+ޗnQ:�61f���m��Z&n�κdW��D�X�*��c.�����l�x���K�w'$���<�1��
u�:�w'9�����P/���5;��X��ݺz����^�ya����VZЧPѥԖhìbf�˺W��i���	�*7�(����t%����(�C�'T��%�i�̮��̎u!��ox���ʔ ���'�k�<k����da�ͷ2��E��)V�rhC[z��JK��n���R����yK�I���#�+.���"��$����'h�R,V�Xo��q� ";�WEl��jT����q�,y�/��������cƵ1��3y�rtAgN�L���}�My�����l�*;c��R�X�eE�Vv�9Rօ��jE��+�+T��q�y�p���lFL'�Eϸ��վ*E:F�J�?��+.��.om}������rv��'Ì1���T��^�����?���3�q���$]� PK�+Փ�  �  PK  ў,J               162.vec�e��A���cwww뵱��l�[�[�l����؊�?�����a��a"�,��"�)C����<RqT�"*镩BU�Q�ԤV��mWG�K=�Ӏ�4�1MR!�f�h�7�-iEk�Жv)��:��Dg�Еnt�Gʢ�]�ދ���/��� ����P�1��dT�����c�x&0�ILf��T9���`&����2��,`!�X��fE�L.g+Y�jְ�u6��6���la+���wȝ�b7{��>�s ��!s���8'8�)Ns����<��%.��qE^�׹�Mnq��y�{�r�)�#��D>��y�K�W�5ox�;��|��)�d)�z�7�;?�B�����)�PK��-c  �  PK  ў,J               163.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=Ç[�&��:�bұ��S�*KoV�6~W�-�� ��+�)y�ٮ^?A�'����S�Z�2o�T��J���ܺc{l��dDU���K;�$N|1}a��-u�Eh�{�_�<��9��ϟ��l�.���bQ�Ƣ\��l���+QJGϝ4:S5!��v�}����׆�FN}R�i�t�'���_�I�/�:�����וי�T���Y��O(�n����x�n���;l��/h�i-�y�c-����yA��h^7�-�^z��l���*zO7���z���ۯ����e5��ڦ����z�:�g��&[�ʾ[�t��:��2�å��>ݲk�l��S�*K�����c�a�+�Y��D��ڔ�ʽeÁ�a�^�j~^��T��H�R�Ƣ��"�x0��#�ȷ�.oip[;�us���ڛ���˄G?���=S��X�C�עr�C�w=u5_��*r
_��%_��މ�m�zƻ�sǴ���w�S��gK�m۱qwv��g���%�1�k]�M��g��H��Ƣ.|����;������+��t�{���v�M�7'�p�ɕ�{4���i
�*Lt;���/��Q½�*ch)��'�?��N������ͷ'�}��<-�3n�w��N���O�gx�q���LSɛ����v��|w\7�Ƣ��x�����k�2���~���W�ط7�?�}/�S1�k�n����/c�ڵ��W&�?CҙI~I�3���|{mϭ0�Be�IE��w��Lx��|�������m��nz�\��k��tH��a+��)�����b���N�e���[zd�߇����S��زSt��љǉy�gϩ=���vEۡ�]�	�����XW�����`�x��~j�Bݏ��/����-���]�+����Ɨ����|i� �Ѕ��f` ��0����_�ľ,�t���� ���)��
�ϩ��U]_t�ķ�*�?����b�ൎ�n��ݡ�?�Y�:"���-%k5]�@G�	�|��ޭ��
m=6�D���Ͽ�O-�:�f=3d^�g�g���ٝ��
T�6�l�q��Y���1�;s�I?w����_�� 3W)��̒@W��.�Lx0��� PKQ ��  �  PK  ў,J               163.vec��ώa���>����ͫ�M۴i��f�M�4�L3�4��u9�ޱ��p~��]WD�������S�2��\ʢ|QA�H%*S��T�:5RD�,���ԡ.��O�(�D�,M��4�9-hI+Z�&��];�=�H':Ӆ�ts��v=����7}�K?�3 �@�A�`��P�1��Lb��h}c�x&0�ILf
S��tf0�Y�fs��|��E,Ίb�\�2�����b5kl��u�g��f���n����Nv��=�e_V��r���(�8�	N�8%Os����<�X(�%y�+\�z���)7�Mn�ܖw��=�� ��|�c��D>��y�K�W�5ox�;��|��)�d)���o�w~d�����PK�a�k  �  PK  ў,J               164.p�y8�i��9̌{7i�#���V"3�rJj�Sȶ9B!�&%�J�FI=�$��am�!��Ù��>�����㟍m����|�����}?���� ��D" B  �5����||>8�@�PH~A���������FAVq�����V��JZ���8#����&;��v���Q(��������V������Hp7�� ��An��['��B�08���u(  
�A�p����� ��󉓎!�0zԔ�He��:	�����(~I)iYU5u��6C�����K������e�׃n�<<�Nx�t��3g�CBυ�\���OH��^���~���zν���>zR�����Y^��ohlz����W�]�v�����������_X\Z^Y�{� �3�����`Pb����w@��X]>1s�X�����H�[T�R�w��8��/�b0�:�����߉E�'������� ��h����ѯ�1�������1��>��Qmv��;L�?$؜�^�i�	0f�X*���"v��M��ʡ���k���%��2�R��ݚ�	Z�KC�%i��ф0)Z�i� (a����L�W��"��úr��^bH���#��T�K��].n�[�l�,�;��P#_�m��1�2�k�	���/��˼;%��$'ڄ��Yc��F�|��-�'����j��G����,��_S�t������E�����s/�"cO�Q����9U��>WUR/}�F��q�ű/
��~ntڶ(�l���ԠZNU��� �����d��R󍩖}��|�cm`�sG�.���ՠ����4��Mˆ;<�����ZOJ��;L�<�.�%|���!�p�O��f���sY���(�r��M��^K��d^�t� lęe��k�-��bV��j����U��pW/���V�r;w,7ǐs(Ë��X���$�k��]G(Y�@�@�[()n�E%w�3���#���Q7b� �0��6�d�UPyG�B��9�Ǡ;�^�y[n��Ƥ�\��pj�C�'���[�ejno�{��"II��O��jN�ZP^2�|���m;_T����i��ѣ���q{��>���*�Ǡ\�����/��+6�Q&�:��k��,��a��NmI�rݮ�a_��=[��y{�T���d)�Q�2���	���#��q>=�N��h�uL�O�g�ٯ�e�Gr����v��aE���h�����@R�.��zj�R���a:'M"`� �W��*v�]��}5i�OD�&Hsd���x��%�L�kx^�x�9��D��[50�>�J+�.�G���;���Py�o�ƞQ�,��|���nϋl���ֈ�i��*�~��ю�#Y�R��e��JX[�-K��}�8z�fwFx�R[Obq×��ڭ�Lɫ�d�M`�������T��B�vn��h�{�#��W�\�nDI�Ph�O6+%��!���Se^w�N���_T���PK
K�  �  PK  ў,J               164.vec���Na��y��������ͦm�4�L3ͦm��WL3�4ԃ���>����s��e���Q�"�e)��(�ET�+R��T�*ըN�QӮ�^�:ԥ�i@C���8�G�)�hNZҊִI�hk�NoO:҉�t�+�R.���=�I/zӇ����� ��� 3��c8#�|��F�c�8�3��Lb2S��4�3���b6s��<泀�,bq��%r)�X�
V��լ�Y+ױ�ld���V�p���v����a/��?�_� �8��r���d�(N�Ӝ��qN����$/s��\��{C���mY��r��)�C�'<��ya�R��5ox�;��6�"��,���U����o��?���?PKg&��g  �  PK  ў,J               165.i��eT���g@���`�!DBB�F����!DJZ��A�����^����~��>g�O{����9�}����*੒��< �  ���"@��������������OHADH@@HMFNBAOb����cd�cgd���q�p��C���@�b�������������J���I��Y�] R\� �� b�{����� �C@�'X�8�x���0���O0���<���<!�"c�Hc�k��0;S&��e�)5������?{NEM������%$�RDT��9y������\WO��������������G/���а��Ȩ��Դ����E�%�e�_�5465�|������?08195=3;7�����������zv~qyu}s{�.  �?��"�ǅ��	���p1<��@��	�M&��c�L�,�K!��_׍�<�4w����Eh���?h�M���E����7�����0IP��S��B[�����ר��"�^�<	<��ZQ����Z�=�u:Ԙ��go3�g�M3���������Õm��.Jp�Ƙ2�>A8?���O�?�&�\��h��v]Er����6�!�ܺ�-�s���v����`���Ϥ���xJ[�QH��*�
���K��41�Qd:��4r݂�rA_n�Ûon�D��%�?~��ƬД&�߅/W�reUQd�������𱐵P4�����o�
X�\T�)�|�f�!�A���F�MB���k�j���
s���0��(��XcJ��N�o�PvF�>���s�9���wa�k��?ىj�5^y��rd;�"	i��mm�̷���Lޕ� �y!xwzhf��m`��dc\Er=�� 
��o��pϜ�s�hɾ���v~O��|s�ku��/t��δ �0�<�/��G�F�S&}�mK\|������v����J3Un9JԀo��hj��&�^�c:\�c5L��?�*�u���z��A1��>���@ߍ~V�vG| ��r�;���ģ�����"�	��a5s��z�#�췃?�Rg���3#�O(q� ��^#mM�V��Mn���/���"z-��k�q���S@h���t�rՌh�xL+�]��5�<:�Xh�+D?�ֶ�x	�3�y��ы���áh�3�o����m����ꖳ�Q�͵|b�J|���͠0��¼�))rV�퍠Mo�|`��_�˙��z�'u�x4�<�b �����(�>�/W�4d8�	�4�M����mÖ͙6��M����~����>;�9p{�.k�3�I��z��{���fz�t��+{�(2����
�&�#ʤ�(4��VoC�8�F�B��4���9�Z��`����C顡 ����� �.ӛ�Q����}O�������<jK��*�#]���k���Y6����)����b��'B�)l�g���"kV��:�o"�>��W���G>�'��m�9z�B�E/p�?�Ϋ8u-cH��D��4�0�I����l!�۵zRt�}�0�j�	����ٓ*yTΊ�V7�#�=$����Rl�Y���Q�9�?�KU�5������U�m��3�#�r�����ao�.�"�,��+ԓ�!s"q�ͭ��܃N�z���R���iA�"��-�
uV��`�T8���|��!����C(�#�I+{��;*��0(��c��x8��KHY�L���)Ij�F��/�wz�w�N��$�:��gtM�CkX�ǡ��];��h��=̜(ئ�C��R�T�ȑ{��o��j7;0�S��:6�J5ʙ�2��F8F�S� ��u�ب�Q�F��a�],8���Α��"ᑟ?ȰIHa�G�0䉉X�i�����͍��vN#n����h�	�L�J���#��#@���2��hx�,���"_E\��Cz�!�G�b�a�ue��t�����^q�^��������-�g%þ�t@�'fL�?��[T،�AvMT���B���զ�]Q{�Th_�g-� \c,���\�Hb��	�h����G�1�zg��OR&����'D�
�Y.o:{h�	�V���6���.˴�_�$�Z0ˬ�d*9F	!��Fƭ�T�%�0t���:K��T�D+��=���l��]�K�+�)j���_�>$��n4�[q �Ϩ/��6���}�p��<6�ί��Yk�?�F
��es[�peEE��ґ��������C�ҢDUbrU�5�E]�f�P�щ�-��lc5����X'`O���Ò��c�"s��bޏҽ�cDG�S�]��ʾ� �HMs���M��k�բ����9ӄ�~9k�%�)�>[����݆MP����L��V����G�A�ϋ��^MX/��ț��a��)>�	&��_��X�OG��}����>�*M��	w4��ߖ��PBoD6�j��_f�:�7�x��g��qn�v3�J�HG�(t~�Xg�r��뾷-�*x?#��`�����_y-s��oI�!5~rF��up �?d��@~7�e�)����YB����R���z)i��Z|�lv�jZ��XX�4�PpR�����M�Pv�3��sYu�	��Ԥ7�����C�ⶰ�A�g�L)Z6�:����m�`@��Z��R�%��ᢸ�~"��e0T�Ct�`A�a���/������?.V�#zytU[ME�*/�l�jL��'w���ON)�[�§g���R"u��ʵ����n�L	ޖE~���#M
�Z�_�	/��@��%��C�/�.~�f1� ��yh����E�呡$Y�;m�6�ҽ���E��-��#�)P�d�8�u�	���Zx.W3��~=;Ȭ rT�Cm*&���%h�F��J/�.˔LB�T��;,ce��1�i�;�r'���.6���l�J>��
�s+WoCۧ\ �n9��@����M���Xa̹ ��\�G��2��	�>��6�?ߥ�/XV���
�^���\��n�}���q�|�{P�s W��RSȭ�̃p2`��A'��
T�C��_����~�g`#�Q��*�x��|d,U�i?שB�D�Z����1�?D}��Eq��i�-���ԑc5BG�6oW�N�i��������רN�>4��
��Eӵ���*������d3,�"�O�"����`�٩n���v�:Iz�t����a���=7�dX_��ԯ4[ޡ&�j4��?C���#����{���~�;�@�C�
s�g�zP�J[�`k�o��)r�In9`v���L��{����=�Wyګ� ��:8u7���cJ��{҉��'����%�NN�՝��+6��{!�н��c�j7Ŭy&��^��8����?�n���|�iF �&#m�|] 	iQaG�l+vo�F f>4�±����"�(�K�?t*�׆1�Wm���j&m��Y�e8.���{n�%�}��y� ��l�k��7�m�d,�a;�-�
�@o�����Xm>��-�zJ�_�V;�p&����3˝en��a�e�5���l�����Q	��P���$"N�T�D��@H]�jTƱ���#��#��$X'_Sx��*���3
5ʝ�*[fD1p��x]�Ak�4�tV0�,����Z@Q����j�c�wȘz�K��_է�e�<W��>V�Q�H���7-5��X:ź�>�+�6/\@�����ǅ<Vv�1����NI��+� bʩ�c�
76V�]���ᷤ[S�Zu�,��7�p�cE}��H�B�M�e���jrC,���E��u�f����e�0|[�R2�'��j�M+:��v�^�{d\S��e�8��^b�C�
��W����5ϯ�}R���;�<���6J��|N�>�\�x��`ۜG�w���TϤԆ�2�Lj�\&��Ԁiށ���O��+ҹ	��N��#'��st�QA$�2@�ާ�����br�J����f�����a����)'������= ]�f��R�otc�_d��í�2�g���ou��{=r�-�.)(s)�% V����De�N�v�M'����ّ�T�a�?���U�*�ܭ��(��ɮ���S�>vFе��j��;�	"I���Ϟs!'���*��{���E���$Hs��髬]�C�ދ�n���q ὂ�	"�A�/E�&@T2&̛(���T^Bt�p4�)H�!#A(�~��l<ٚ���Flϡ;��;K��/�	M�����n���!o���UT�õ3�>3�ȡT
�tT�'��B|�G�iZ��Mr`�qtjŮ� 2c����1�u�?hZhY���O�1�2&·�� �c�2�s2(yOc/�%)��d�%zy_���,4�!�!�/�0�P�3*�+��Ә�(i=�7� �� �w�e��BZf��������'p6h��Z�en��2�P����>%�Se�x���&��ֱ�x3Ĩ���I��j�#@o� �NcQ�g"����=F�#0~��5��;s }{���5�Tb���Η1dJ��p���\~�Nl��rK2ą�Im�@L�FAS51�FI�+����hm֫����+m>̈́��):g�6.��ę�s��3���$�A�BC�Of�Z�	��5���d�I&�Ց��m10�5�=1�RP�q�����bu�c54sB��KeH	c��1�|L�+�GZz����K�Pk:"8	��\��ŋ9�&j}����e��*R���l�+�:�׳	�;Iԍ]�_���r����S:>�n��c��&����5�5K�"��<�A1���/�j�n�,W��T�+/4����B���oè�Y��)mi^�F'HU�Ih �����YS�x&��!��OSRrC>�:
?h3hy��17{���c��"+��&�� !0�����O�9�������p_�J�v�h�^��X���:��2�=9�Z�\�H�q�kh�t~�i=�i���.Mi��)y	�5��e�"$���9`���fo7i��|Hn鏍Q�	�uCG���5~(��`ve<qR�UDw�]�h$�M>������m����� e_�|
��f�t�B�Ko�xt����&l�?x�7:���}�®H;�u�q�U9��;����`�)(d�U&p�$���{�l�J���
�Ȼ(��9��G��s3vep�
؈S�I��iÑ��lN��smý��c3I�H��e��%�=�`�7��	${*��F>S���A���� 7|�:�P2_�υd:��k�*j<b���w����9/W�+*o�����;��k��ӈ:�_*Aj��O�«S�͡�]v!��U���Yߐ9����>7|5��)[7Q��Կ��h��M+��;���f�]��������C���b�9��*�׶�^ϣ�3?�\M�q����{�G�s`�P.,'�嗆<�JF@'�3�d�4[�n6(���Q*��'���.K�ޘ7'��4���?/���q-<>��Jg�b�������m��c����@J�"l=���G�9��b}꽳&^,�da�
����S���G��	罉���k�+s�̓�@rH�&po���*e����I�y8�N5t&s;i.
iH4�lЧy㴢�z��	X�IR��.�>\ojsǭ"���l����3��I��*�s� ���z�⨛rؘ����y�ׄ��pi��w�8�x�8��>��ql����fcFY/����ص���Y���G�_����D���a��+��N�-��#  �n�����(='�}�4�tpm_����i�-Vo�"1b��"X�*�ơ�KF�Bu�:.Q�+�/v�i99�K�ٲ�=�0o�<;�D�V��z��江���$��筜�@��3��,1�B��:3���@�C;�-����8:e�)�vW�֬_�c���;Ɏ�_d��
��Z�%�M�\��d��,�L�Z�=etWL�~�����U���s#��*�޳L�jQ/�C.m`��V|�f���'87���g.j&��)g>�-/)D�#�d �R���mx#�]�q��w(eN�-��Q�!ZO[jV#3'b��G ��)��y��*y�,mY�͡���o���[�菦27��R[�����nLd2;tDꢌ+����c��H(�𚬽�M�ơ��aWA܂?���.���l�vl0��]�r�� �
bq���Z�����:r��F���{�i��{u;%�_S*���s� Lz_� �gpT<GPk�8jA���#���r�PQů&V8�I��[��z��;7!�"�*[�n��q*����l\�i�w��Մ��� Q;]d��:�m����<�LQyUk-vH݋��[���_��jT\�	#��0������W \���req�8��ٖ:��.j�h�/���&6��7��s�3�j]ӁۀrCr��?���m"^L	U���`��jea�P����d��${�5�֨upK\ߒ����>���+�ᢪ.o���O]��mϙ��tW��,ڏ�,A��s��[�F���~}�i��a��i��T�r	Ht~ ���W�Ј��[?��E���v����?韊�sp+܈ű(4�eʻ'�U%:R�2�Dk�|GZ��t�}�4��p��F>���Pc��^�*��$R璃����s.m�Z��i5�:i�+i!�Ȑ��B��Ů�k
E|=$<j��6�99����~�P��.�W�H*J8�_�?3�z����M��B�5�ϓ�.NA�k͋0�+^�Y��u]�"������/�ǜ��'x��z
7����y�z�$� ��_�V�����9�j�裺*���׳�ؖ���%�c��J!�S�����tt�{:F)��6Q���<�|�^s�S�44|��~T�����)ŋ��O��]'��Ҍ���PК����?#�~dς��E}�J�<��w
��c.�y��9`����/�q�^%׬n�TMJ�b��{�/=%)��֐pt{ܨ�5vh��^*i_��V�ÃR��lm�c��:��Ӷi^5��>V��K&MٮW��V׵��P���oS���+�o���4�Y�e�^C�7�椯5�d�5r�?Ǭ Xd�Uf �h��� �C��]ކ3J�ֳ�:F�-\>�E܌�c浧Ĉ�*1|&�%-���s����!��lSe��Ǐ����u�]a����9_�ʂn۹���ZsJ!S�tU��Ɋ�߮e�B�Lq�'7�u|A���*J9�����Jv��y��������x@G��Nj|#�L�� ����e�)
Sɻ�F5Ѿ�X�c^�gȾ��Q�~�M7��)����#c�U7+��k�vBN�+�u��u��W�XCidX1��!����C���X�s��6����^N�V�fT:G��B?qԸ�&F�Ž'R��kJ>Ͽ�g?��xwy�O���-���x�F�O��e���U��Xw�(�֎�Ji_U�beo�\��d9�j��*g��xmgpp{uٹ��iҘL��Lz1�wEQ�Q���Ŭyx�����u�����7�n�$[���/?�Ĩ�\>�5N��������F�~������l�z���B?/�g����sp��x�#�Xi�U'Ę̞�>�`��S��̌�����Ti�|�v+u���̵#yh74�2ƛ�K��f��ƛ?Gs턎���r�# �
��f� �ڜ��L<<mu�¥��ZZ�^;��V���{q*���%�6;S��9š9S�
bB��D}��p���W��'&�O�Qe��=�����~꒩?J��1��$��J�=5��6L`3��YO�L�ma�
Hl�۠[��!�e9�̂��Ű��c@�ȗ�q*� ���{�o[�~)��%3��_	P��2vѨi�+2�Kԍ��\���k������=�;�Ӑ��U��2���K�B1��Q&�E��eʰLI¸y�s�|�L"jƬ�9x�c�9K�}q�k�?������D?�ԯ�̹�Bl8�fzeη�-�WoEH�k%���w*rp�����	�Ň+j*�(��Ǖ�(C��_x�EG�����#a��o9�-�K�`c�`���=ÄE땜��G�'R��:㖣�)��2o�t;WFt�5Ϫ�Ʌ�i6Sk@�Ҋ�����_MCosJ8O���b����ז8�ݏ��Q�[��b%��2��1�C̞<$��h��k\j�]�9�ݔsL�H-/���`O2�1�3�,�)����ޖ��RV�!豳�Ų;|�%	9�����\�|4��
^}�ᾫ�ԅs���T�)rN�����9�D�>��J)�/*�x��/PK/'!B�   J!  PK  ў,J               166.pՓy8�y����)�;��5�� �L�%���4���FO��br46[[&�hQ�#�L��I�i#�J9�r����j��}��|��_���y�����u�z���� �  @���H$
�@�P(-!IX-�j����,AI������������*e��"�X��A�J��4M���o�1��/1��*I���D}E�\� ���!P��A�� I�N�\��� 8�Bc$V�/�� A08�@����q���*z�5�>(Փ��t�Z˂Z���j�a	ٯ�r���d�uTC#cӍV۬ml���qu����������?t:8$<"2�Bt31)������4΍��3��sn����WTޯ�>�=����iG糮���~������щɩ�w�gf?|\�����/������.��=���3���U��h�%+�������>F����O}b	m������ٟ`q�I�́�|2�����,�n�e����/e����vz����+R�N~���v�N«�3��-/�Эtpa���n��Yh�$_����
w�)_7j0��O��F��K7ޒ�M�{�ql�����ǚ��Nnr;9/\�ƭitc��1?ɰ#���t
�<��Qz�!��H-�Z�P�S�5�0������gk��l���J��ܖ��a�9J�~O��'؄7��:��푮�5��d;%Sg_W��Q�Кo������kUٺ�~(�{��5�p`=cP��#i"�^*@%>�k�'٘d!6��%�� �x��FwK,NM���k�Kս4�<a��l����2�~p�+����e�uɾb�9ٟ5�wW�Eva���ʨF|�<W^4���R�1��k+�@�)���Ľq)%�s��>eג2���:���Wn���OS�NVj� �l0�P��n;���L��`�,��d�DGލ�@���+T.L�|=��/ڈ5��u������r�r�ݜ��"������~y��c=%�>��-U�cy}�@h�ر2���wvď�219�������}X�Y�N���a����J2�ߙ�a4j}��F!ż�����|�H�D�Y����S= ���T�j촟�ދWj�q�'���4���fd��[��Q�s���������!��[�㽲�mA�n���xU�#�74���u�7��0�s��\A����R~W/�D2���\��9p���#-*�� ��ɱ=�����u�ސ�VxUuW������
ǧ�~T�ٽ��]�^�<G���ұ��4���rN�8`�ل���#���z���o4����YŅg�ҳ����zo�*�����K<��@�l��|��c_��~&�	�Q���bR.��+!7�h	��Fj�Z쫳���5���E�!�f:݌S9�: ��۟��r��7�S�y��	J"�屳�Y)2���Q�P�u��ŋ��r�'�P;ƌq�����|�����9Y���I۬���_��J�"F��>W�SZ�D��jX�q�������|�zc5�n���uS�i�I��\���!�\�9��CW��mT�Z�(
*�=a��u�����PK�rC  ,	  PK  ў,J               166.vec�g�NQ����轌�K�n�.�%��D'�Q]�Kt��`0��^KnV�����{ND�����
T$G%*S��)�jYDu�5�E!��C]ꥈ�Y.�iDc�Дf4�E�GK�Vz�iC[�ўt��d�Y�BW�ѝ���m�Ⱦ��?� 3���Ӈ3�bF2�ьal�������$&3��Lc:3��,f3���c>X�"���,cyV+�JV��5�e���n6�Mlf[��vv��f�,a7��a/���r���(�8�	Nr*��<�Y�q�\�R>���r����oo�[ܶ�#�r��^��0��|�����%�l^�7���w���|��)>g)�d���������~�R�PKzXnd  �  PK  ў,J               167.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=Ç[�&��:e,��a�QU��Վ��?G
����w��(;���)����=��������nA��U���\��+�����"�t��+�}b�$89g����/c�L:���0�X��?�vݍ���?]O�%�i}����^���
jν��P�Tӟ=g��yyR�����*�)�=�G��;f�ת,�9��g/[H�v�N��'8,�e-:�u�K��a+���-ۥW�u��M�v����>ݔ?����ۯ�����[��]�{/��������>�(�u�p�ܭ��~:�����,��Ң�u�����_ږ�n�d�������+�<�~AjF�]�EWх�B�=q��蘬l����?�e��-�Ԡ������Jox����I�W��<��豤-�"ui5h,�b��_�q_έ뺨��P�r��9���v~7�Q1���w�c	��y���9f�D��+���h��v	�!d�=�:BwN�.q�qj�ku-,�����Y/�8�mV��(�z����X�GVJ�G�ex�8�;Lt������)��s1�H�S�=�������זə�>se�U)����>��l����[zf�Y1����v�'��M��~j�X�[��%5�X
j��?�f����}E��9fͪ��fԥ�_Be;ޥkwx��[������1_e/��&���#���Y�
��y��T����r[~�>�.��Ek�6�$����O-�ս����Yӊؗ��v���]O�s��NwY�;V�L�M7��^��p�䮐��Փ]ENqi,j���L3���+���xk����]�{�ޕ���,=�+e���LC[�s.�>��n�9�Zx�F.�������uA�F�.<�3Ll2��J8Q��K��]Ԣ.	��x0���V/�l��:���uo��ó���r�j�9�mz��3�&�_�?���7�RW���`�*�d�w,��1��"��z�]ў��'U�j�gg���7�gWقi+����[�S�N�˸��:�
��8��r�����P��&<��'�z��Y6��j��)?c����w��~�Tm�s{����[9;Xj9�	]�R�ðyw��^ՏF�ii,��H���xS��R��{*��ʓw�����Y�kޅ{'����SA��9ǥ��:�wLdx�eS���W����i+��r�mvO���7IMZ�H`H ��� PK�bծT  ;	  PK  ў,J               167.vec�e�VQ�玾vww���������86�`�`+�؊�`�zu�K.��?l8\ΉȲ��P���De�P5eQ-���נ&��M�R��)�A���z#ӄ�4�9-h���ʮ�ކ���=�H':�u��w�����'��M�����@1�!����#�(F3���c|��&ꓘ��2���`&����2��,`!�XLKX�2���+�*V����c=��n��&6���lc;;�i�K�f%�e�9�Aq�#��9�INq:_g�Y�q�\�����"�r��^�y3�-y�;6we)����\<��y�S�����k�����=��'�l>G�/Y�������GV?��/�wJ� PK�M*ed  �  PK  ў,J               168.pՕ{4�i���3f\&RL���ĸ$i�!J5d�t����T;���)�m71˄"wf��f��H�D��҄u)�����?�v��=g��|�z����|�����n@���� a  * � � �B��4��b�pD<NY����J�#���#��Σ��303�Յl��[XYY��9,�\fN���ib�X�2N�׶��;����6@���@64 `N �@_1'��o��$
��*)+
*� ��p$�PdY�<�  ��[�@i0��D�N�Щ����4D�F$b�4��u�A�&V�6�K�:��]�V�{x���f��F� fpȷ�C�"�EE���?p�H��G�S�i�32��p����<����²�ʪ��Ow�
�ꅢ����-OZ۞�w���x)}������/#�c��?LL�p� �=������!pz������(�t@���e����)��R��H�MJ����3h���X�"��O� ��	 ꀸ��D���Y�AIL'�ur9�����P�柫�+�W\�����S�%�jD�e���9��Lv��f.�粹Nl(�J��Ѱ�!i�3B��-UN�I���}��ʂ	���m���K�n������I�*���3���qR%e��mHH V}�z@�,<:8Ĭ9�9�*�>e���,�b/k:��2����6��[�9�!k6?<��H8����C�woM��bȃ��͹.&��)�zr?��
Nܵ�������!i�?��yHys�u�"hOj�_s��è���9ut�/|Ed��t�K���*H�T�Y�J7�7�^j�Iq�C�����g��,A����o�d̮��ȐȆ
.�M�aό7y��HǼ�-��|L@�O�DuQ6�����au7RqK�6�$IKo�N�;�胃�l`6,�ɗl�o��|V�$��D��J\�_��g�s��_� !E�e1���zbLm_���Uǆ����2#�suaLh�#5aX��~̔��֋�������(7�l�]���ةТ�o�w�`�a�{j7],z��g�$����Ѭ��V�?����Y[�)�{^����eIR�l�x�|A`e�o�uA��].&6}�;��<�ᖶ����4NC��KƻU_���m���h�����1m;�����m$�.h�X�q�^�X�&^����� �-��o8s��ԖC֯"�i��v�R�4a��7S\ݨq�$��^��u�6��Ӻq}6f�F�ռ
2բɘ}cW��Q���ck��\JC�e��Э��dY��L=c���S�ˑ�m�D�ϭrJ���7!�+�F/&9��_�eg�����|/։�-�(�8��j6)����N��8s�D8U�`>%X�91�k{ad+8��us���r-�+f�ܱ>gX8{4u���3�����5.���%[����!� ��X�G�4E�t�:�Y|��eW�׎�["|�W��thڐ�xqy�d�.�I^޹�F��UTñ=[��A<iI��&Յ��{����ro.\���L'zC_{��6�&��$�l��ة���.n�FfQ�Զ�k7Hj����������t��,���RB�ޅ9 ��u���C��k�6b�[�^��t�k����WPKf䤅b  @	  PK  ў,J               168.vec�e�VQ����kw;vw`�ݝ`�؊5*��-؂�؊=b+����������܈,����B��Q��T�rʢJQU�FujP�ZԦuSD��(��hH#SL��,�y��zKZњ6����`�Ѯ�ޙ.t���AOz���}�K	��� 2(�l7D�0�3���b4cҟk7N�&2��La*Ә�f2���a.�����,a)�ܱ\�`%�X�ֲ���f���&6S������e���.v����c?8�!s���8'8ɩ|y��g8�9�yy��\��㲼�U��~]�H�qS���y�{��S.��<�)�x��xi�J��oy�{>�O6�#ŗ�_�����G�7~�_�N�PKB�8*e  �  PK  ў,J               169.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=Ç[�&��:e,��%5Uyjrx�[�]K<����L>��tJ޾�E��6~]뙧<#�v�����4?W0T�����̒˛�^,�ZHoG˪�:�b_��@^�y��1��������~P����i6�����߳��xl��A�ho�g���;�2�����l.lo����~v��ܘyQ���,M�U�Sa���W�褉�"�!��"�0{��(W�5��v5w�Y��ܙ"����ޯ��m�e�����.-�o��|���j���r8qn��	{-��g�`^a����Ҏ��m_�s׬ssH�������.���\�pa��e�����WIܯ�/����B����z����,%��������Nså9|�Mo(�XԵ �� l/������������ٚ��}7�^1��wfk�:�y�ϩ�Y;���������@���4�.S��R�����J���dO�i��Y������w�yv1���t?���-����u�E��IgE�D���ҹ�'���嬯������z�Ǣ�������V<I�� ��~�ߌhAٛo��.+Z��62� �$�P�]{�n9?���z��Rv�J�K;s�g��,t��3��W�z��Q��2�E]80s��N��?E�.-fH�=�.���G�3�_SϞ�ml������6���9�N7:�M_|��=Ὡ3����dPQ����ʯ�w��n�{vNՓ�2����V�y(3Oz�{\�������y�+�����I��QS��&�W_��b��j�3�'���n�i�J��3Ev�<%���L�8�zYM}��JխM�6�<)2��e����sW����q�t��:����ο'l���������X�+��2���s�
�<׉ᓹ��G7�⻮,�'�^~T���f���:�3�1�"Ӏ^@�ܽ�O�\�#(�]ûC�@�����9_�V�����=��[dw�i����g,*~�n��9>KU��.�-qO� ��L�����R��:r�;q_t��gQ�h���m������WN�vqRɞk�Lz�9��_M��|�cj�~�r˥�f�� ��J��ޞ���ϭO������������k�&�7�a�q�`OJ]h��<ыo��艹f�[��*��߬x�U{O��:��5��i��3	�c��n�f���@W<���M PK:GF  +	  PK  ў,J               169.vec���A��w�ںv�����-؂-�b+��-؂�؊�؊��]w|dx8�Á��e���(Gy�T�"���������W�:5(�&��M�Q7�G=�>hH#ӄ�4K�hn�B/�%�hM�Ҏ���`�Q�Dg�Еnt�=mz����/��� 2(��`�!�P�Q�pF0�Q���1vc�q�g��d�0�iLg3��l�0�y�gY�b�����rV��U�fkY�E����&6���lc{V;�Nv��=�e�9�Aq�#��9�INJ�<�Y����.r�P���
W��un�\ܔ��msG���y�Ô�G�1Ox�3�󂗼�y-��w����g�/��k.ŷ�o|��3+�_�7R�PK�b�Zc  �  PK  ў,J               170.i��eT����t7� 1� �JCHKwJI�t
CH
C�C�tII� ��H��t��֍7�Ž�{^��ڟ��:{��8�� U�U��� ��� i �����������������--7�sN--�k6N^0����n~��\����GH@""�1�2��?� �E� r0О�dhdh�= �_�Xh�-����C=)����������������`�a�3�JbS���<w����ŅH�tQiL3���?y
�~������]@��k!a�2�r�
��Z�:�z����ml���=<��}|C>���GDF%$&%����g��~+*.)�^[W������gwϯ޾���ɩ�ٹ�����ͭ��ݽ�ӳ�˫���� ����#�?.tLLL��p��{�ǁ���\R�̅�9_.�T|nM�_���u�	��������7��X������\� !ڿ�a�P�XДO�V��#`�)��(��Ȭ�6���?��-�Y�6@�PI�_#H��lD)v�x A�i1�/�:L�8ߺ�e�*4$���v�#h��z?d�C�/��uW��ł�B�b�z��G��F�ϐ�ć����VW�yS�;�&a�|lY0����x[�p�ƾͭ�c��E�z\���'W��->&����W<������=R���nb��k8�����x�:z�:�0߻a�-Ė���7�TB�n��%|b8Av�I�Z�^���3��O�Z��Cݾm˒�Ҕ�}g������.��)�Z�5��i��D#�u�����^ͺq�+�ţp�+��� #�/޻����{�.�RX0�jcP�h�;��t�YtTX�:痔T9Y�4%��X���W���נ�,�m)��[H ���w�=-J�ӟ��?92��^�t�����F��=����W8T��\���}TT��yU5�K�,�os
�L�O��ot;ײ�ތ���
Id�9+��qr¸���-XPxa�\x���yVzu�y����z<��*����?�����~�X7G�i��x��kշ^�'X���K��v��y����=���q�B��&kaa�����nzYXkϔM^��%=]�u��p���$��1�ͮʪ�ӈ>�䏚�m����1cO!�9A��iV��u��LƉ��!m��@�kW��ZX�Oễ��/R��������G�m����k�fcR&���YG��S?Ҿ�-9���M.?�d��4�G���B��6�t�g�C}�l���;��K�k���ub�L�A-iU�F�2�i�k��6�rL	K��];�a�%�m�4�|��#�ә�(��g'$�V�����)��D��Ev�J�Jߑ�!ԉ��C��4I��#���G�n0e"8��0�%c�KkVu��e"O�,w���YF�1��aY{�qd�9���H�G @z}	)� ����$�P���U���1Ǝ8��Pl=�d"��������|���K�n����":�}R{����9����*��i��yk��T#��Tz�o��[W��7N�P�sl�a�k:&-��.8�E�'���nvfb�M�ō��F�1�������0���i,x�%Խ�Y_ڰ[��F����0�Ύ˵ۭ�~�Z�>��w��%��O����G ���Kɗ��&��;M����ʭ�|�|Y��ך�G�Z�A��aXq�<�}���E/���E�m�K�5�������eV}U|qG�xس���9)O�������S�4����&x������`(D=քD͆'���Z)//n��-�4��K�ص�-��3��n��͚6�-%��D_����*�c�q��H�+��7*�n_��[>�f�sL��o�'��p^{i�˹R�����DW�}��#61��?dK�E6�GI%)����1�F������=UN��	���cˠ$�/N ����=@�<Qe���D�cx�"�LS��)*�Os�v#ÛI��ꗝB�M����{3
����̓��3+[�XLD������~b�)�`����p�C��j_o�9ɔ�w�e�u*���MֲI�4���T����iqZ�ۼ$6y��g��xo�<�x�ʴ�,��"N�@4Or�%�@{.4l1�
�|�����j�7b� ��U���C��D�̂�m��ZR��3r�4����g��/�;�Q�\n�����'��5�_���A���N����G�l-n
�����E������^��h��(��KZn����l���#f�&��7\1ټ����As�n�a��68������]�c8rZsf�WE�2y!o@�W���=�o��{Q�	�it��6�&��;/ͨ����Q�=y�R�d��P�h���ENj�!�Q=�s��=�W�je��K��z�.P
��zx"U\���=n�$��ܝ_�@�&#�����,>���4����9��pR��"�	$�;�/��h�[2�f_��[������t�C�zu'3�>���=���kr�v�m��-ګ��R�H�$ƛ��\��ɍo�	����+�8�������ьD�'�*�?��,D%i
ް�$��٣+Er95�����!��[O�2?C�F�M
���*݉�Q����W<��;��]ߌ�҅�y����'�+	$�r,��7kY��A����:��.��J��M*+dٳ_�dbO?Ұ��-��<�z��kP��\�,2��wO��؋�<x�������`�����m�.P߷�G{�E�����N"�GB2�@��k�\V�u�ίA5�w�����Y��1��՚S�N�p��R�j16-��T/#�7��L�K��6'?Ѕ�p!�9ͪŧp��t�&�b�;�{�wu^ϖ�*З��K1�󒻐���k2-Gf����УEά=\�!��2SPnV�?Bhi.Y:��LO�}��d��M��B�!�6�\�Go�؉�p^�i3n�!�J�r7���gq�u��LÐ��
�҂d�l�sm�X{�*:�w���t<��N�S[w���ZA.���F����&�k��]�؃���p�����?E���I�q,���AMj_X�m:�\�����q��"�QF3o�fgry뢺	+F,՟�j���eo�W�����ґ�5��5k��NG�X}�P��'���x/Ϲ�xZp�����Ҭ��jkʭX�EE,�)[���6�(k�tW��B�h�Hdh`�V���ZҴ>�wX6{������Đy'J�"z�$��"���M��q�i~��=��.%s`�ؕ�%G�T�ɵ�N����ȧ��jf�'wr�'�=ô({�f�;��~7 ����S��o�$!�4���U�HNJ-1���@a	��b@�l��pN0�S�=t0��/�M��ղJ}�ڭw����TNy�!��:��~#�e:Cc��H.��z���׮�����+e�ּ�����E�L�Br�MFQ�/ط������˺�j�"<�v�� m�����w�	:9��E����%�ă	�1�b�͛�ъO��5~&��yH(/T����6�/�i�W�&��li���to������D��1�R*�L@VTP���h9�qV����~�+���	�av��(��_��>BFB�c�`ڒ����t�	y����њo��`+���Zk���C��I�d�b_� ��y�"��� q4h��.Aʬ��p��$hԋb�m�G�Ox 6TM�zb<-�\]�����)�� L����Ɉ�l���g G��qLtڦ�߂�[D�w�µ��?��gkzx�6�FN@d�j �y�[re��W�Z�+�D��ḣ)\�zl_�$c~<�����<
[�:�]ؠ��[��m�۠�o� !���0~�oY�b�Q�w�$��O僳�<&�_�x$��<�7�)��
ͣ<���9��2&�j>�ָr��bDW�Ë́]�AuԛW�K�r�@i��|嚡�w�,��݀32t��<�#�o_��<��8�1�m	=���?��4����b�]���C�%��OE?�Gm8����qxH��I	� y5b��a�7�1�x<��;�=^�א��Θݳa�)A �(ֿS0�If�Y�HR)4��ŝ�rK��x�����$�6�+,����L?=�L(Q	�P�9/�k�ey�J�A̋�pPz�.lSR�Zi�{�Ul#So��ie;�;�h��}xǻ�Z�f$$1���q$N��F�M�����"߶����I����OjZ̀(���� ���Wl y�4�+n�B�[�0X>�D�dL�\��Z\��`n���fx�m���(W�ž�d������
�"ԩ/��w�}P�
iy�����]��c��V�ϺC��bO����Fm����^@@>$�A�$��b���ֳLg���d}Q*T�2ҿ��4�}��d@<��jۗqc�̎x���R>"�FV�&��������7�#�1���9KLp6��r���DM˙7�����#��l���b�ˤ��P�ΑԪ���Uj֤j΄���4_�솜�q�]�8=ǌ��{Hֹ��m�9	#i<����NĮ�;���ρ$~�`^��?��R�=3.8Lv)�݉�R��V��(����qn���y�\�&_�"׊�Ȫ��ԇq+.J#
�Y��e�(~j�Ď��������p��j�.R&�t;r�B?vY&��*��LI���Yz��/N@�`�:�W�[�Ŕ�jޛ��y��#�k�2���(�)��E� ��˷n	�V�q|�L���U8ɾV��~&q�e�,�_�V-�k� U�S=$��r�ރ7�R�t.��&i�F�zdSr���, ��ݰv�����z[�,iφ��kG�6�z���	�w��3{�a�6 ����U͚�~��C��>=x���q��n4��p�I͛�
�*��U�dNf�X���mp��v�� �󧣒>�HC�I
Y�l�b�����ȇ�X�_���R���s#�mE:�?݉7A��:-�;�O	�9|3�:.e��"^V�ҍP�ȕ����6�)�lRh�]�����Y�j���G�q�
��7�ȥ�C�0��O�����B�=��o'�~5�0��6I�+�� �`��(nFdd�/��1%'i�����tf�#<D�@M��ZI�19��#�t�V��Qu��'�=e�z�5�����Hݲ��_4�^r��;;��-�i�*;D-(x7��[u0����1��t̄lH�Iv��Њ5��q�����0��A{�����mi��c��׷��.���iZ�F}!J�9�5d���)�J$����[���i!\����dw�����%�w%V}aw��ƿ����\q����8��������Ɨ cDM9�ҏ3�o	��>x��?�g�������HS��).�/r��*J�ٓ�T�L�H`Dge�"�s0ZB�Y��rމ�ex@��R�ʒ�o�X)���%�&�;��J�����f2x^�`˽�xA���v£�G
/3�v��Ɖ���
�����VI���uk����wN�Δ9��6.J8vS�֛C"s�?�|sػS���꾯�B���?o��oJ���Uݠ�p�a&l7�`��������q
*Qz�x��acW�(�oJ]E�����Gl�wq���Z}n�|�@���́���n�#�]ɞ��3���2}�g��<c9��[�����F��� �:�
1����r����ɏ k�������+��0Ϝl����[P!�VM���n2Eq��d�
����B Wz���y/�oj�[m?�!&rJk��C���Y�������v��G��e���.VH���WN(Cy����(�E�T�x���N&��[��-(*�X�G��C׍���/ܝe����i��tE=y_��w6֘T,2$����ԣJt��ņ,��.ϩT��U���<O�����㾪�'c7���m~Oa,��\v�>�k�P@W`���N�����RM��}�%x����"�'���lQ�{��2��F��o�u5(�x�ļr��^��/���'"��Z�{(>Cش�jK�C��D��.2�cw`��x��I#�/;�����,U���ɂyc��LK�����V�=�^Q7�u�?�Ÿ+��1�Rj�:bQ���$����5eUKrr�N��$sJ@���#�S�_tB�c�%��.���e�,%�,#~5�+�\��Z<R�Y��ӞS�Eg�_�:@��ƿѴ�5���vQ�`mhAK��j�g:T�is�
�A���o����ϭ�� �*�5ӿf:��C�i��i!�0&�>aΎϬ-Kq0׹g8Z�
:�뙢���r�������4��s�O��A�UT�R��fr3�1�	�`�[:��O֥dw?��g_���e��,ܻ���*t|�j!\F]T�LV�<���/H� �$E�&6H�&�d�4�ʖ�XJ�#lTή������
��P߻i��.��D_����|�d�<�-z�h���(�Q'����ٕ�Te#pw�P�e���yQؔ�K��E}�i䣔r����#˰oly�<G,;L�5�I�c�E��x���\=Ԫ�я@����J-(��������k�A�^�>���0��y4����d1��:؜M\��ۇFa9
�
��D���w�'E:�A7,9�Eu��M��=j�/@՝(Z�6<��0�5j�aʐ8Y߇� �Vs:�=A�r��$���I�,��K�'�9���L�*>�BgD:����ϼ���_8�Z�ྛǕ�Ћ���q��w��]�e�6�֜��,����x�3u'c<�.\�~]c����9��%hp)B�#���ʤ(�*�}G��6()C��SD�Z��W7N�|���S��E~��o\�H*��M_��3�h2.2��m��v��N�b��ǔ�f�V��B6*�6xbtx�"��^��
2�)��h$F�
Tq��92d5�CG؝#��J�b����N�4�tq�Ǉ[^�n���cH�Qg��F��|+d�VoJr��������M�e��Kg�.:FJ�L����4�����+hϻ��P�{�$|C�3Cf����f�	#�GŊ�Ű�	�?�V���,��~(����0����)7����=� �TnN�R�Sq�����.@��b�S_�7��34E�(E�{Vt�BmK|�W%w��ui#5��w�����e�PV@L��&7^<3(j�e_�[t]��Z5���^�\a�h�Q}�đ��O������Gl{XD�PQu������Em7��]q5���K�cD��S%�0�5����?.3'wWB�d���K�&�j������7�Z��u�2����p�v3>�����~왖ʼS���a�L�_�r
� ����o�]�ݮ���M\ݐ�~m��)�4m�Unϥ���5"�1ע�J�,C��4��,ŻV��p������WE~e�'S���^*wV!�.������V(������6��T�y9no�Ə���
X�E��$��,Z?����g�BW��"�G j��튜V�*Sd��AJ�0pY�o����r>l��W�q�}+��G�L��ӁDM��)�	�Ю� �O�>�),�0�G�$/1.��z�*w�^�D�6�}ʾ���tҜF̌P.s�9}����t(�{��/w�/���Bt�ń�T/�<��$�VJp��'��~e8�7�d����Rx%��N�w�%��jb�A��A����(I7�����Un0��_h����8=jI	l>��$i�vQ����	g����6R����U,�X�P�ݎyA�I��dUtv9�N;�B��Cw�왯�S${���^�
%�#):O{����_i�<��SXɼ���b�d��/o�m�C�^�z�L':m�[a�R���[��&d�S�$<��4E�{q�s�wel�s�/��}'Y�~��ih@/�ZV̈́�;֮��ü�}=���30�M((�����V"B|LR��u0b@��;�db$��W�z�y�:�^Ezl�Iٴ�T����م:Ǘ���U�"_('|�w�������'�Y@H]�bc����ġng���~c�v���=u=L��t��;��̋b��z��B���OI(�T^ׅ��̉F��TGK��$Ha����\���O6j?���_�H
t� K�k�,	��,��ls,���T��f�=����#��|c���������j�!uӾ�y���P��.��llr�
��PK�Y   �   PK  ў,J               171.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=Ç[�&��:e,�{R�c���n��L��]�<w�g&�q'7^���4f��=�nZo]����d,T=?.S�Ĳ8���E]I\�艭rC�OR�]�԰���_�2u�=���iV�8�i��1Gݳ����_[Ĝ����[k�4�<�;F�p���_����;�����h�ՒGa�;-���2�
�,ٽ�ILq�����g�]��*�E]�0�Ə�W�^=��rf�ї�3���[=��7�6���s�P�j����3ȵ�n� ���O��,��^{]'�=��c���u'��3�h����Ɂ��n9H������ST�#W�6�&e�G���O?β�=y��4�D�������)m_�g�ٰ\!y�
�k;V2x'�:�4���j��.�.�1"/�=u��;�ӓ��^)#s�2�F�7,����s�,�<���7�?�S'�Ι��ώ�9N?�K]Y[	$NY��ǭ�FI=���W1�T�>�U�<{ꕛ��@��{�K��-N/��;Iy�Ո�ƙ��,oQ��u���u�Jc������/����1{~�<W��`�S�ce��/c�Vx\I����g���jUOU3��Xf�/돭�>b���C�Z��f�?�쥮_�[o��i-3�5QbG�F|啽Z�]�3�і��W�{����3,�<z1�����_ֻ^�����q�,(Z�����볶��ui�U�@�x�����y��=�g�J�<f3'L6+[�s�=-�3��0\�+�Ȼu�3?���Z9�����?�Ù�޲���%	�-6m?��y����t>_��h����"x0�͊�[&�<�.�8�\�?у���1����N����Z�s��4:��?�����ӓ�!	4YCcQ>��tkp�
c�I�S�Ze�65�o��n��y�ד_�MV�-�����Y!q�CK�?0�y�����!��7o:��7��j}�!us���>}�������[v�j�z�����e�������+��x̣�����󳞚����z+z����3fԨZi,���*���G/��zy˴O�6��+>�ܢ���y����|O����U��.�3����Kt���=�u��D��ŏ���B29�5֜cc��:�����ӏ�X-�DL��� PK�KҬ  	  PK  ў,J               171.vec����3w��������-�b+�b+k����b+�����?j\�G.���LD���_�
�S��T�r�D��0���Q�Ԥ��C�,��]}w҈�4�)�h���"�GKw+Zӆ���=��;�uvw�+��N=�I/��ڇ���?� g�1�n�{�)f#�h�x��v����D&1�)Leә�Lf1�9�e^������,b1KX�2�'�BW��լa-�Xφ�<6�&6���lc���CKlv�.v����c��=�!s����'�$�8��Q�g8�9�s��\���^�*׸΍,7����qG�r��<��#}�����%�l^��R�;����~�O6�#�/�,������Ώ�o��_�βPK/I2�j  �  PK  ў,J               172.pՔkX�U���]plL��PBC	t��u
q��!�4C�L��
�Q`!R��&P�5�K\��{r�._���/���}:�����=G��< 8>l ! ��h��j��Fc�(������8==����hiF~����������ƁbaA]i�܉N����4��3�6w��bqz8}}���5����u�w��l �xH���<QЫ ����(4F���]P�   F a
���~��H<����M�F`l�DZFn���r���	[��V�����l�b;���ˊ����kX>�k�?����A��xQ�1;v��Jܗ�?�@Jj懇?:������N|~2�T~�����s�KJ�*�\�����k�75s�歖֮o�v��*������0���ɩ�UϞ�̾�� ���z!�H����s�H���ȋ���lh:D���ˍX��	�ȄN]�-}p���+�7�+�?����8��O0�G�䠈�w�ϐ��Ӯ���g��*]]m��[}�Z�Q�f ���O���]�l���!��"n�/@�T���XR�f�}�r������s޻��!�C@���K[�ݵv}�g9Y��l%�%-�Tɡ�p�^�a�i�������VY���d�G+.�GL��L��[�URK��wWG\�HcW���p>6&�1n�[�=���#Dh9S{%TZ�Y�cF�6S�]r��ߥبySD�`��6�f"�^GR�jHQ:+a �.�nB��Ҁ�B�'����0Yu^�V����}�����;2F�A�}'%���S"�����}߼U�⿞�Wd2ҫg�*V�����!���]f�����5r�Qp���%e�D}�s���o�����di\.�pn�#�dN��|�� �y�"ɸ�m���b�n��T�J$B�@H#�� �ݪ�(�F�Ɲ���~b�FÓ�eb�]�]���,�4*�(G�ÏcfFN2T���g����%B*��x�`úxMр����=5aD/iYG���s��㞷z��f��ի�ݦ��A�O&ү_vaٗ������kj�|X�9h\����z*^C��*�<={�H]����m9_�ċE�3ᲈ�5@�C�ie�u�d�yP��:g�\�x��*�W�K:�2�^��T�{��-��:��I8�m��/���ꒋ��h�&Y1;Ǆ�;Rn��%R�K3*�)P�%���R�ŧ����K�����m'������Tۅƈf4�>;�o�ݞ���7>�׾�<�8l������M���Ę92�K*��_��'����s���!z���c�A[!�������ü�����@��N���S�P�d'>�c`�.�6Ïw�>� ��VZ�w������&7(�����[�4xv�&�t)�Cv�~�be���w� 6̃�U��8��o����
J����:�was<}�Bn|}��&|;�+:h#����t�O��S���t���ŵ�E�1�"葺�xzq�K���k9��q;K��[L�zk�����ȫ>�'p��9�(���G�282]V�X��P&诏t#(4`��� �q8Q�vkZ}m�c���ƴ+��x^��F����tڮ�I�A���<FCͽ_PK��N�P  2	  PK  ў,J               172.vec�e�a��=���������
�؊�؊�`�`+�b+�b돚s|\2,����q"���<�(��7e)Gy*�,*�UrW�
U�FujP�Z)��]w]�Q�4��i��hj��ݜ���iC[ڥB�����H':Ӆ�t�;=lzj/zӇ���?�Jb��`��2��`$�m3F�2��L`"����2���`&��͜�(��<泀�,b1KX�b�.g+Y�jְ�uYI��ld���V��=+���]�f{��~p�C�G9�qNp�Sy��g9�y.p�K�_�+\嚿��H�qSoq�4�;z�{��m�c��g<�/ye�Z��w����g�/��k!ŷ,�������/�͟��PK1AT�`  �  PK  ў,J               173.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=Ç[�&��:e,�8U�ܽ�aΓk�o�����^��U9+9'��݂{�g��s�rLf���S�;$�ՀKcQ5�y��g��|�<�����5W��b/�l�f�w���uY�+U��6T`<��K��@WєV>�ۘ��f�1��\l����^�޽`���MZ;?�=xPt���:��m���E^`�-���)�BƟ���3퐞�m���\��};�*S�9)=a�W{���x�_Oꦸ�n�u	��X�ŀ���2O�ʑI+�>���g����Ƙ4�ݏz����<S�):]�����y�y�>%�M�ק�u�ƴ.�U��4�a�%����If��{p�p��y�s�g?ʵ���\ܭ��S�y��e�]�3c~Ϛ���^0	h�D���x�b����iO4�u�N^fi��[��{�ʣ��bwo��9�m[�I�혜�������N�[S*賀���ݓ�m����׬P�[t��"����^�q�^�w�{�F���_�z�+�fD�Sz*��*����?����]��T��9�����m�\��Ni�Bgg/��me@��b��s\ʭ��K�����'��`'s���_u���ݮ��Vm�ź��m���y\]�9��n�]���'x�8wjwѹ'�����=��K�_����K���G>>�ޡ ����u�ON����W�P�Ƶ�ka�	7��0V�y�"�_^��w�i�	��?�gީ�z=_-T�}ݫ{�%o���%������ds⾳����,i�ԥ��	涺{d���+��n��cO�<1Rt��}���M+���/uz���뀲f�.ז�g:Oҗiw����\�8�+�b��+Zgg���z8��dᆛy@c	�H꣈E�f�kZ߹^��u���	�)�Q_��z���T�Jw}2_�gT[u}.���"�w�����/PA��WSᗳ��Y0�����LC�N�(���ө~��'瞝{�L;Ow����%��?2⿶��W3{[g�/���:�N���!dͻ-�"s����v��I~�ſ�6=�u"��QBq����S��?yi遲�'�;m���nx�u]���g�/�=��~��K�]?4�XԕJ�4��ky�[�P�1�u�������gx����b֗����3���ޠ�J&q7�.��3�}�����z�e�Q3u�;�X�s�ݢe�Bj��ǀe�+!{��� PK�=�'^  =	  PK  ў,J               173.vec���Oq����^_��WwL�+�ٴi��f�M۴M3�4�L�G}];{�����s"�,�?9�(G��T�"�R��|TqW��)�5�E픢�]]w=�Ӏ�4�1Mh�
�̮������iC[ڥ\�����H':Ӆ�t�;=lzj/zӇ���?��� ���!��ag#e3Z�0�q�g��d�0�iLg3���,st.�����,Ɋb�.c9+X�*V�����:]�6���la+۲�خ;��.v����c?8�!s���8'8Y(�)=��r��\����2W�꯹��S>n�Mn����.��������<�)�x�^ڼ�׼�-�x�>���s��������;?���S�;�PKjm b  �  PK  ў,J               174.pՓiT�W��/{�j � �!��"�V�Q4P���5H�
��,��b��U+	e����("��ܠj ��� �DP�������=ﯙ{�<w�uɤ�2���= B  �@�� �$�B"�h4JA	���������	�������@��56��6�!(��L�t:�d`ekI�16���h���^YO#ȴ�F �����6 ��P(kH�>��� ~��HZAQ^P���P(��a0y6N�`�*�����Cj�ai��Q:v�M8׎�������r��
=}�*C���������L{��Y[�����������;�v���&"2*:��IGxG��'��srO~',�����������U�5��._����z㧛m�?��P��-���ex������WSӯg��.p� �#��#��`Pr��D.``p2�����SӦBa��+��:��/p��u]z����{��K�Wd���%���|xP� ^H(´>�4�,�k�V��qD� �J�?�2��z�ҫ�SXi�0�|������銹;��g�":�c3�p,{�!�˒�i�g�(ܡ��/��(��y 5�pv��UkH��o?=�s�-`m���+iF�H<Qx��%�k�����\m������'߫��PL��ݛ��F7i�Ð�v�9��L�Ex�C����YF�4t�&�VLz��S�#�*����
�ԋ�8ɽQN>%��]SeI-�1�+�Ğ��VfXv7�YϹ#���P�3���=yRégFq�����Y��Ӎx��;���v�D�n�Sey��V��t�;��o�팛����������b1�u�~{a�CY�5���Ta����-F����1�%>η�\F7��j�nf䊈��<�d�ϓ�է���Fdk�[א�C+Lu���$^�R2�.�	����kDK\t�ڿiҒ^C�㉧�K�}��]5�N�2w��W��y������m݋v�n���M�|
����&+w_�6�hܽ�~I���c�ډ$�ةw�)͒�l_�=A#�s&n`�0�5�|�̈́/�����RFg�!�=�B�S$�,:�j>�=��K���I��Z���
J+�=��"��o��w��l��n1�uk4��E�EC[,7��af��U���A ���n�Ɨ 
�GU闏=�"zĺ��u�*�&��fRPT�ԯfG�����'^I��k!�l陼�9g�u��9X�##����Օ���Ե��L�����y��)�o�ו=�?〈������<6�Z����W���Ͻ��U�L,�����
�y��抃��� 1�N��_��_��f�R�l�d��:v]��|����'��:�:EB��mb{R�}H�����u�3��/��,	("($��lj:R�bc�}z'	6���C<���_��'�Qu?���Q�����^���&d��������}�v��µ�fά��Z��̴���#&b�)�*7�~��;9>��3KD��!5퇑�t��1L�s=7��o�^��=�)eQ�iN�����`0�z��)䜯M�k�6��� []�~��X�&��<�Pخ�T=�[Ձ�-q���G&�A��&�S�^������V޼SZ�4�o���/�Q��<��n�p�Ӹ��ּGy���h�>�R��ʺPK���  a	  PK  ў,J               174.vec�e�Tq���?�kwwwcw�-�b+�b+��-؊�؊�؊�jv�x����0�漙�Tɓ#O�)Gy*P1KQ)売�
U�FujP�Z�β��{u���O҈�4�iV�fv��-hI+Zӆ���}��vݝ�L�ҍ����M/�M�ҏ�` ���l7�=�ag#�h�0�q�g��d�0�iLg3��l�\��y�gY�b��4�2]�
V��լa-�R�����lb3[��6���ء;��n���}�� 9T���(�����'9U(�i=�Y�y^/d�����lsE�r����fV��6w�
qW�q���P�<�'<��y�K^��捾����G>�/6_#�o)��?�?������oV�PKk�9i  �  PK  ў,J               175.i��g4���G�D�Nt�3���{	Q��.��D�%��&:I��5z�N0���n�r?�{����u���׳�~\x\<SQPV �� hO���bc�`c��������RҐ��P0�212���3��s2����s���a��	I����4<<<BBj""j��/����� �E�a�� �I�0H�{LO��B�o����10��qp��	�����00�11��01�n�����Xd/�ɵ-qX<(��R�qY_û)u&�؄�<���S�вsprq󈈊��Kȿy��������o`hdlb��������������c@DdTţظ��̬�Ϲ%_K��+*���5465���������������_����������px~qy��w}s�� ����E�ą������.4t���bb��&��Ʊ� g
åx�Z��c�9���ħb�`?����߁����/��͵ �@{*) 8C�J�J�;�|��h�C�jt�\y����A���lɷ��.,�X�G�3��兰L�����T�C)��+��!�*�5�9�drc�D�ګ9B��7g��3��B�R)�����[�թ��|�b�vٷ��oa�6[MD�	�B-�Q�@� Ӷ��������3�r������Y׹�yh�����k�3���"�3t�F~�-����1��� fܮ��y�c�Z��>�'�
5j��h�0`MI`T���M��
0s�� ݥ.�D�Tf�D4�:�?L���g�%��@,(Z�	L`�1#�2�V��
�媲��F�����QO��9}�I��1�g�u��⢐aы���L*S���尥,Df����˗Jɘ�e,�1⺿�� �$���%��Q�eԡo��]9j�/N�YKy7 ��J"�ލ�zkm�F�Z��S�FǤ�~�5�G�r��WH�Յ�Si��A/��PՒh�÷��d)�7��<�&�$o:y8[[X���%S���!�FkH����Z�!k�����BQ�Φ;��=�43���>wq&o$�Y��Oa������,4Q�8{K�����zI={5����]��.���-g���MKu"��ۡ�d��-����/*���z�ǘ��+�˚���˦�(�C�u���j���~A�����u�R�.�iE5"=(ԫ�Z�v�^s��0Q��y�uk�;ڹ� @�*���s�p��y��u�ҟ�)��b�A���C������5v�`ω�:�L�-�����1�K��7���oñ�C��԰�*�Z�.*=�vH6��QҠ�q	��=�#`�Jd�H�8�WL�`�|T��1�����FQ���e�z)�m�E��b\3��B@]�Y�}�i�5Ilv� �Q1�&q�ܶtI=k��]p���<w��+Q���������}�il'��{Z�tV����&�D�g�.��l�4�����RH����/�+Au�ۈ��xS	��Ɵ
l�����Vv������1���^c���(��m`x���GJx�{�v�Z?LCd� ���RJ�l�Cg�F$V3T�t�ή���aW�])�92?w[O�RN�䍾t�[�'+�6N��9N3	^SN�G��Y�p]������c}�����X��9��|��"� �(��y�`�灆Xg�/YF����X��HLR��H	L���$7~ט�{jx��R��\'x������1�S:���Ύ���S*(W>t2�g���]XD�*o�1�֎$�jZE��F�J�}�W#���Z`�낪S9
��R������/��c��{�Y��bDrȂ�������\.Ų.SK���P/���٤�L�m�Aߟ�qFD�H���rU�M�i�B��~�CDL��%�G2�ZX[�MW�.\����۶���k��J���^l�&���`W5�tE�0%��Og�(q;�|���y�5=��g֑��)�"*��k:����^�6/#S=�*E�ɍ����ю���noPl �x)r���>b�D���@9a���o۴�������<��`����|��x���6Ī�.�XJ�z[��e����ߴc�Z�{���\c�U�Bl.���u��
:����Ӂ�o���(�h�
���MwVrSo�Fƅή(A���$�HT��lI ���
�8�����I�W�;UV����W����?
{=ل�?.�g��������*��x�
��KZ���J_l�ލ,)n�y�`���G-�`�����:��r�Π�v��\��(4C�1Ձ�A-���r��vNԱ�YBꖓ��p��$�@-X�X���rj��z��P�l|�%߲���C1}�*`���﷽A�˲@I"�b'�7r�fi�����=Lh-℥��m_�|Wb�Q�T��Y:l�L���5��<C[�aك�[��f\�n�+����7~�8]I����Q��(H����R�9K��]����T��'�A��K�L}�����J5-��lO��_j���¹��lM_�k`�/%�!O��-G�\�列�ʈ�D�}����t$d�✏;,�vJfdwUk�ϖ$*a�=�)QM�R��ّ�[�*�nk�`�g(?{[�+d�ӏ�Gj9�Q��c"�#_{��l��v�Pi�����j��� c�T;��w�3�Q�4�W�s�&��+n�1��N�MI�+a��4�-�w� '���S����!�S4�/�eA��]'� �>��n��,}l�K��=U�y��tC5/���䉮�v �^�܉٤[jE��(�-�����&�ިs�9&�Y�&�Y�-|D~0y�E�����p��jt:=��yɮ"$�Ѝ"e������1"	��)��$-0mbjC���6��?�sb�����#�gx�# �_U���d��YÀ���7	��o�ɑs�#��G�ߕІ��Ҏ��9�jFlh�!+rɗƇ�/�:j�����D����}��l�ٰ�B]W�mw��m~��w)��ep�"����W*_C�h=o������u>�ض�%%~�9��zO\��[�h�NuR߈�li9Mo��ZcQ�{�[�6����sEiPT8�{ ���ϟ�qˁ��&�0�9�]�����{ߪ�޴��׷��s�޹�v'�%cx��'�
�ޭS>�d���k�B�� g�XyK����F��5���N�s��y�'����a ����4Wdڛ�f�R��~�����]�A�f��U����U1�J�d�y�K�y#q��u�ć`6����)�M�W�$ė���+�6E�7=��k� ��=f��X�)���N�-����)ꌲ��{�.�W���4&�4����u�R���~�QD��I0A@B�z���}篼���a���Q�ݬ�:J=����[)��x^�\�U�İOg��<k�]�׈�^F-J��>d��Io�_�����r;��
�J���C�Ц�z@[��ݚ�\�0��Ere���7�����2�h�[z/�g��v5Y��Fm�l�� Vۜ��,/{�噠�4?I1������ܜ��4k�vL��e����eZ+s4&�������!�g[�71���ŷ�ޅ���;Z���@%��t+L:�1�A�����_�t-h�'�·��0��Py�&��7�����(c1F���7l�l�z���@��a-e�2�Nﮣ�N�?����!r�w�����X�-�}��>�� ���Y`1Q��xV.~���9�իLO" ~@��~�&ˋ�q�嘷}`�r��?�����<��������I�"���Ƭk<��U{�L%��Gz���h��RCPd�ʱ�&�:����������@�a����~�����Ot��4<a9[u�֚�ד,w5o��rlJQ��8�=(D��"��5:#ʍA��c\��A���*� ��򏕅���<| ��p������am���쇕F����}d�3��Ĳ���0�l���A�^	g���a5�O�(�mt��Q�=��!M+G��r5=/PW^C9�(�+��)ݑq��_����t��KEң���� <ņ!��X�޺�|	�mHV"�x����Dk�?U�e֥�f�r��9�+y�K��9s��P��d\�ΆG7e�M�W��x�e+Ɍ~��אz�������/�� q�~ϫV�G�@5���y�1��>���P�:#�����KlS��o��z��/�o�'��J�]�f����,�9	��$���}7TC�A��>C��ޥ�C�Hlb{�ǖ��M4DlwA�0��/Y(d��S>I�R
z��ԏ��-z&LM��Ce��l6�H�F�\q�]P��<�ހn�V�oPMjs��T���y��9z����[g��K)xqh�+�ڳ���}�Մ��Ǌ���+ ��#�B����;�}-��kg�E�~�8�jY��bz�����ߪ��@�Djh3d5^.�陹�v��Rof�g?}�Ye�=K��1n� 訒(�4�{>�C1Aݧ��!�`M>j�l�*�.���;�I�&_1W����k���1�Mx�r+8G����k-77�����^�K5�N�=)�6�M�'4�����	��8{�t<�γ��	�F`.E�ip�
����c��j{����k/4����(���xv�ߖpޑ�|���[	���ə�gM�@��N�B���l	���ϫ2'����i���O!�
��v�Rv�f��5K���xX1?�uL��8f�s�3�i"C�x��a+�P�fC{f�^���,hp�$U3#������]�:~�F�&���.?�j����%��u���%"��-
��NHM`��y���S��b�YP���s�v���U܍D
�lk�s4h1P(�ƶ���Ne�&�F�<}B:J���V7ly��������k2b�������k&�A�ɽ*����b���q�/.0��IV�T���֪����� �c:p~ph����Y@�y��[�H��4�	�o��#�Kԯҩ�c���\y����r'y,�'x����xQ�����`w��`��H��թ]�!&镔�]���n�X���K�<��Vn���	]�v2������d�J�2�b�|!�5a���4�|�-w�R��-�#��0D%~3W�N��1Wi�M�n� �W�s	'�"i@�CF�o�,!������u�t�n������eFd�0�
Q=븐���h�BH��;3�h�,��W��ط7�11p3�f��pmUt��P�`wgt�3��q~��&i�p�([P���!j�meiȗ-@R���x�}*i��̓��:�$�pQ	�yc|�@�R�Y�Y�+ϭ�mO��?^�ʁ�R�������p����z�6��!K��1M�f���{��?V���9��8xWͻ��/TVS��EqJyS��z��Syp�/&�_�l�Tx���q;��͒AF~h��:xP��g�����l���E��P
�a�e������vϛq�9�a.3ڶ�+��S|�&a"�������U)ޞ�u���G@�W���D;�8�ѧM�㷆5U���9���yudB�w��_�����������7�>ޗ�\e�yZ�k<$���s�)Y���7�T�*��A�B�BCd�a�g��=�W�������*�w�l�#Swf8���>3ι��)h�� �K$�T{��[S��[��H���o�I�+͹�U�(*��1f���}�)w���E:V,�%@�k������h��WĒX��m�.��?�P����1�k�-S=ߵ�.8�o&Z5�V|��!���,�9yd�A_~.އI�z��F3P�s6 �O�S�Uw�U��(G°�5����Z���Y�=6bh�:���F�!���E������@.-Mp(���y�̎h$���_������SբDA�>��#�t,=�ʪi_^�z@Kvq�ͭ�e�YQ�ʮ�)���+|)y�P�گ��Tm�33�ؤ=�
�Ͽ>���G=��j�D���4(l�
v���F`�)EYej���;]����i��:��-BL��#Sza����S��	����f�(�9c��8	�N�p[�hh�@ߖu(Vu�ww�LU�I5��,��$����D5�y6�5��3ȶWt]�b�����D�)�8p�jt,��Q��|RN>��k5�F>�o��̅�͟�%��|���i��d�i�kJG?�����O���5�J�;R��J\���/f,���	���=}�� �↿Vu��,����}
�=�6��I�V+�������1W�I<�,�j�;�3)�򓚊�xӜ�69�8����c�Bb,���.~T�74�lHJ�o����ꏧ�;9�+0Fr`��y�f�`�4����Ͱȧ��j�&ْv�<�ǳ"��L.��?��u4��uSj�f��YK]= #�X!�"�ל�q�3|Ӆ;MQ>?ަ�5�K�����=%�vLhϴ� ���Z�cCH��+8�ϧ��0G�Q��/=��4\��--J⸨u۷�+H�7N������Z��A|�wL��Wq�����#Gθ
&U��s��=��)co��rc`��|�D)>:�w)t��2�w�G�7�:K��}���}��@%�?��&m$߻�ώ���{�g�k6�9�H���a��.=�|c�	|O�4*L�@��d�xm���1h��ݠOhCt�4 �3ԫ�+^��2�r4Taj��R�3,���⏀#CJ���Z/�k���M�q��~��J�u+y:�,����'�퀑?��V�����?t���7���B`��~X��󤨧C��ԅ�k++~�!6@���L,i�r��Z,��N_̪��!wG�V���V������୳�?'����{-�V��9~Y~��������N�g���s�0�is���G�aϴP�Y��d���"ӆ�!�] ��S�7�YN퓗+�Lj��>�j@�/+�9�$���w�z#>�;����MG��D��)��A5=o���#�QI�W��O�q_Đ�"��>�Do8��Lfn_�Wc�i|@�Z�i�0}��7h���tw;3���c�#��{�^��^����,h��:l۞��w�Ю�?����d����hɂ2�r.J�%�{J�\%q nū�2
4�.Ik+�6���O?����z*ntT���[��.n��L#�>�e3��9�t�vH2���6�.�\��TL���+s����� ���`��G!�#k�������
��3���`�w��Js0p� V^��$��N��@�<���Ǡ�E:��5�T[Z_����	���][�g���w�	�T��)���Eƞ���k�"~e(�{,%�� �`���2�癌��V��6X�/�c]������ٚI����B�5�ca$����>�HD闼7ju��� 3�i��1�5]N>����J� r
�b�l�#���n'e�Y��_/���ӕH��N�X(�;*c�3�SXo��Qxy3c�vԍp�Y��њ���'��Վ��`ʸa��3D�<��5����Z�B��`mU��|˕��h�zh�\�%�V4�A�|iz�-�^�\����xKˁ�R����h�V�-��������N�/�I��,�bH.�Dʛq���9���qY�P�z��%��n���S܌�%���6��FcV�I&�L���;�F����װ�=S������Q�3�����5��M����@�ep�`�T��%|��#�K<�;O7��G���n8�y%��
�.�|8��C���Q�#۪;6�o�L ��}I��gA����RWV%�|N��ERNԣ�U1cb� �F�s���/Pm�W�)��:��K8�#*c�F��C~B���_�O$�<-��_!_����
t�}z~���D�7��zVt���-������Y1"e�sϨ����;+����W$�k1RG/�g�}�?љFhr�qE�{�0�s���_h��u�[��/f���	o�φ
\��.}R������1/̵��G�`��2��!ו�8L��h}!r�M�kw6�q"7��xr5@�$cQ� �1Anڌ�JH��@-9~�c��20����c�J�}J�V ��z��"cF��]��q��#�@�0�L(����ڑ	ҁ`�A����+�N��L�}M�Hc�����A/�^�z_��8:�4�x���q${�J�8�-���PKnQ�   �   PK  ў,J               176.p���/7O7F&F d�������������������G�����GRH�_DVJ^NVJFFAEO]AIGYFF�\S�����D^�����F���d#'''7�/���������AF�̌JL��̂���0����P�����������T�U������������([�g`dR4tdLdW*1j���C�i�AѠ�T����8���%$�T��54�LL��-,��]\��=<��CB��#"��SR��32��KJ��+*��[Z��;:�&M�2u��3g-Z�d��+V�ڴy��m�w��u��ǎ�8y���+W�]�q���G��<}����W?}�����?������X�%�3;�_�L� �,���lB��쉅�JF�"Nn<ȩl�A4��"����CՏ ��}F�ǚ���c�b�afF� �=Ç[�&4ui,`�p��6b��6U�s�-Ы�z��*Ҵ�-ȪնV{��Hn��	7����k=�T��R������"aї�U��C��u�׳�~	i_���l���99r���<�+}���W]BzW�Z�H�.��E]���ҝ�]M�Z�e�g����m��~]�����5��šr?=���� ���}[n,�{5-2V��L`��qW���G�07Ґݿ���\򸭁��u{M�@�wKy�_��X�E�ޔ��P�2M���]��?��j�����.jOԼ�;�~���[q��H��U���b����:�ò�yz���x`��������b~/�e�c�w�}W�6K�gM�g�Y�j.�_[Z�(�1�Kcâ.|�y���)a�{V5J&:�`���ovo���7��?�\���y͑EM�/7i��e���^z�SWP���EW�S\��a+}�;�z���lv����=y���v�v헸}��K����Z�5\W�_q9Zh{*0{Mtt	`ăَw.���z�MSDC�e+C�Գ���^�������î��b;m�x��u���&�S�y�y>�� bfd����CuL�[�x��a��-���ߺ����m�ڊ>�����ݯ���&�/����nX�=�U�q�I`'��ޏF���y�*F�9b��G���-�^�S���G�IZ���y�	�E��/�=�v�c�3M�wj�m}�W�=m����ms�+&���|���L�Y��I�!�U�f���tפA$obJ�<I���֬{D��� ������.�z�p��n�sB�*1���T�/�����=��'�3>�K}�`_��p}q�)���?'�cv��i�Y�?����s�t^�/�0u��,�EM�
L�eF�qn"�G6r�}h�����[�����R�8q��I�Y���7�L�����_ kAդ։/����Lޜ1C��:SD]��r)���7�ʟ�4:w���O�r�/-��R��rh��܂��%�K�j	�V��VepH��?���G�ʴ�mw7�8�g���FN"0#dc~��\�n.C�	7_x�� ?5��#�i��#�ܵ/3��c��8�NϮ�gf����)��1z��3\�/�l79WY�S��R�/e���O�|�ʷ��U$X�Pj� PK֐�v4   	  PK  ў,J               176.vec�e�UQ��������:v؂-�b+�b+؂�؊9��؊�?�:n�<��a�?lND����QD�)K9�S!eQ1���W�
U�FujP�Z�4j���^�zԧiDc��B4�k�7�-iEk�Жv)��:��Dg�Еnt��]O�b���C_�џLb��`}C�pF0�Q�fc�x&0�ILf
S��tf0�Y�Ίb���<泀�,b1K�\,��X�
V��լa�7_'׳��lb3[�ʶ�4���d���^���,dqH�G9�qNp�P�S�4g8�9�{��"�l.�+\�׹��qS��6w��=J������y�S����y%_󆷼�=��'�ϑ�K>��|!����������_���PK"q��g  �  PK  ў,J               177.p�k4�i�����gƐɤ�0ƨ�2�a˥�m�c�m��k��U����%&��[�!�*4���2II;.�ʤ��5;:�ۛM��z���z��<��s�?��nN�N  P� � �@�P
�� �Acqe��Nc��2��&YG[�D��7���SI$����Z32��ޚ񕩹cq����pDee"�B�0�u�o x4h�A= ��xP��9����(G Q�UR��
�@8��#���7N� ���3����N`$��Tǋ7WxvO���;����$jh�ZM�ZX���f�l��rrvqu�v��7�g�w�A�;w���y *:���#�)GS�xǳsN���/�))-+�8[y���r}C㕦�ֶ[����=����?~��xxdt���K���w��3���^  �����+�`-z����x�b�Z������1��G~�ś����
�}�Xu}��$�j���ء�d���'�� *�쀩N� I���Oh�T���UW4ǐj�c�N�w<��H�$O�^J��3�h�ħ.�Jq�%��tC�	��4����Ѥ�C�I��HU�ke޴|��6��<\׸�7s:��MW��=����<Y>?��ek<:��D���Ȥ>�-F�� ����JZ=ֶ2˽2��e:~��H^�Qr�4CZ��j[�n�Q��Z��b�w��ƣ|ۯK擿�ސ~�Kͯ�@}9Vd{��ёG/�}��6=�9zz1[_���〺������
Oj2U�6�e�p7�3
�&�b��^�.H\
�gx�X��iu'@C�j��x-7g�>�VbZv2�����M�[�=�iV��rl�΃�nY"�Ǭ"a�yNuc�O��3C��,D����3���Za��I�(���*�5�e�-h76/-�MM>S�.��c�����H���D�i�z@`GJ��~��z�@������ɯ��mo4C��W���e_�$[g1"qņƪ	-��=)�ht٬���5#��}WUl���w���a�b���/q䶞ͫγ�f��?%�f��65k���1�B}3��t�8&5�cȧ���WC$r }��o3j*4�&�M�8��ߊ��MO"~���ؽ�5u�	98�t���\�0#�z������%�n[fb�{��K��d}_y�0#����Y����A�s�%��ER �'�#m� L��p:*�~��6!:��h�����/o[��]�U�Q������8�ͨ�nAH�`KY��x�����)�Dr���si�Z>�Π�X�𴫳VJ�aƗOU�·�v��oVܖ�%����wE�O�c�F��Q��"���k�	�ot|�g�+���.��f�rHs��,�'�����IJ[~TDC&��I|ou�{X�w0�(l�Rn��rN?]-�H0�Ad
�R`Z�A�a7��~��	��F�*��fɷ����M+�R_xA_ZH[xD҅��:�Vi���)ԉ���Ή���}(��''ޑH�I�z�7�R�r&r).�yhl�5_�s�/�{��B�7�şX㪦|,�G��/uay����RU��31��n����s�)?��+`^{�gP|��S�#�������A(_ִ���|��V�L	�D3p��l��"|��U���PK��Ȓg  L	  PK  ў,J               177.vec��kWQ �s�Z�k���;f7؂���؊�`�`+37�)��Vl���x|�����snI�9�AJMjQ�:1	u�4����O҈�4�i���5�[P@!E���i��֮�ޞt���B1]c.t����'��M�ҏ��7�n�>�����c8#�o��(}4c�8�3��Lb2S��4�3��̢�2f3���c>�\X(��%,e�Y�J��J�fkY�z6x��r��f���lc;;�i�K�f{��~p�C�G�\8&�s����4g8�e�<�.r���\^��5y�ܤ�ʘ�[�6w��=�S��<��y�S������|����|�#�l>���1|M��M�Ώ�o�������PK�#��g  �  PK  ў,J               178.p͔iT�g��/{ a�%&��	��@���Tť��E9� �*
���A�
cPЀ��A�PV��%��Cܒ	���g���1g�{�_����Ϲ����S�0�/� !  ���(����H$����0��#c,�z9��z���
[g�
��ʊ�tpZMsuu%PܽXtOgW��% ���c���D+"�?�m ��!$ŁZ)@н~
�� !P�D���uu� �B!0(��Y�< ����4�17I���
ϣȾ�f��.��K|rZ����b��=��ҕ��d�{�]��[��%$4,<"2���u��;w��MMK�ط?�/y���������KΜ](��x���r��u�7nJ�ܕޓ�[�v�����?0�����ظbbr��kՌ������w^  ����yA`0(��B�
p08��0��"���$�!޷�Mv	V��'w�ں>�{��������������C u̓� 6�l��N��\��G��N�G��X���-r�m?�Y ����n�J'��I\S��n�M߁�q�����s9x�ص�Re��2�]��	��*�3�b�汚-�~����T�h_2p���$��8�}��9����zԽ��@Y��-��t����擲&�4aC冕��Ӗ�t��r��3��j�{Ǿ����8x��>G���k&�x�;,���4�wo,������)E�����<^��\�9�|����5��O��e�H�l�<vE2S�Ař��9�IV�G#:R�0��<���o����W@B>ò�ئ������p�%�fӢ����^��%��L�@�����I�PŏsU���'E�Utp1<��m�}���r��$K�{��f�	F���7(�_�bF/��W��e6p�����K5�a�[�ɡ�x<P��+�Yu`��6�]���c���@~ڄ_>��[�P��xW�r���REg�8���" ��K�_O7,�� ��bJ_#ay�bW�d����=�_=w�!�=:7+>���E޸`��deMN+J�*
�y
� ��d(���1���t�K��S$����b~�F����Fa�!��R�}4u�6���r2����Ot�� #-�5���F��`��q�j/�;��qӐ>�b�3M��+-����Z����q���_F���m-��{�˗��D��߷<��V�b].c����Ҙ�/�܍B��
|�zi������_k��u��d�{�0~��y�v�*ʸ�?A�����۸��54n�YqK=C�2HK����T�h�F�x٪v�\;u7S��ĥ����2-*����3���f�ļ:7TԽq�Ǌ�2`E}{U�M���H���78����-�K,`\�1�ڵ4f=/�5�b�r�i����>���c��!�^ۇƋ�X#��u�bݫ"���'�faL���zC�#�A���2~lf�9+����/℟���c������%��4�Kj(���'yȴ����5��y8�U�K�ܚ��(��1ωE��F�AMpv��s-tm&I�fq"�.ED�k�������w�.P����_|��y;��<�^N��i���&��rL8K}��i]-�����ta�uu��VJ�q��:rȖ�9rv�ƽfO@�M=�1�(��mӝ�3��i��r��	�rLdZ8?�W�/5$�ӒB�z�"��X��? PK`a��  �	  PK  ў,J               178.vec�e�VQ����������l�[�l�l�vs�Vl��u���b����p"�$��ET"�2U�J�<��IQ�5�I-jS��ԣ~�E�$��z#SB)MhJ3�۵�k���5mhK;�Ӂ�6�dg�Еnt�=��n����}�G0�AfH�'��Ӈ3���b4c�8�3��Lb2S��4�3���b6s�˼������,a)�X��Wȕ�b5kX�:ֳ�f���f���mlg;��n���}�� 9��,�<�1�s����t��y�s��.ȋy!.��\��*�q�ܤ,O�\��6w��=�S�����y�S����y%_󆷼�=��'�ϑǗ4��i����H��O��;��PK�Ia  �  PK  ў,J               179.p͔iT�g����ND���E�@YN@DhD	E%`�"�@i$��A@"���uБ�aT(ApP�9��E@[�jhE*�@zf�?S��s���u��}�}�Pl���� P �h�~	�PG!�H4���6`���F�zqxc��xcSSs������Ԕ��lG�:::������莴�&4���n�`H�0���ǡntP�@!��:P�n�4��C~	���08�Bc�4�� (�0��4�M���u-�=V�2GK�,BY�?�x��@�<!Dc�`hdlmC$��8:9ou��˓����7p�gA�>�b9},����$��ӂs_��_�(�de�|��+�RYqIi����k���ݭo�����qۓ����޾���/^+�GF��'ި�z?3;7�����@�?�_z�h��0C�yA���܂���`!#�,i�(���"�C�=��~�g��k��5�_��=1�e���o^/ ,����N��Opk��#z��9��Tĭ]l�J,2bO�QhŞؔ_����� L�s��S�����I�O�1q�Ip,&�䤠� �������.UG?e�n @X��?鬸�FO>�qifNY_<��̚�`:��"Om�t��C���O�.����Sw�NuK�9V�cm���*�(F1���m�Iv员T������y��y�bp{�˜�
�|*��v��4)��������&h�3U�{5	�@ttr<{�^�S�
D-ۺ�mL�m_�=���z~��"+ɇ�z[fĤJ4�$;�{��>(z3.�ٝ�.'��#nT��6��П�4���$l���iV���W�ce�a|�L��,I&��3�q��=�q�ø���j��N5v�"S������>���	�ǹ��CK����h�c�'�����˦2�0�H��"�e��ؽ4�Vap��MԳ�b��u(�Y&y��}��2����L��D��0�[����h�����7�Ѽ)���FJ���v�\�����|	�c��l�qO~�ǐ��غ.ӆ~�V��a���w�ٷ6��*����,3|�f-�y���fw�^r�P5�Ť�7��na1��j	�B�W%�7*U��N[�.�O�uU�͵ĂKAȎ�����/�	�i������ᴕ�H�6��\�y�m�|s�[�G�pQ�9ݵ�ǻA,t�b-�K�YHT��Ou�lI񚷑����-P�By�4^9l�ޒ��(��VV�q|�'4��&QS���[Rv��ki���]9�N!�G��H/�d�S�r�䅒}�sVc��	�\�����c��&C5L�?E&&� VM���5O����M��Z�ksL�m�N҇*[n�ћ����\����5m�YL��W�*��
n�e��f��	�w��/Jwy,�*��+UaK�����W/PgFV8
�H�w�&�g���	��#$~�Mmn�]��KK{N�o�@^Ml��w�G~r���$��)w�{�� ��{Y�j ��=5�`���c�;\��c��鬑�j�7X�+*$���Yj E:��}ܼQB�y��X�o�\H�޷s�٢�X�v�f�/?�y��-9uƛjV?���Ǩ���I+��e-N�aQ�:0�`��E.��4)$��"�2���3� C��l_�Q�׀��k�d|��u՗#���Qc���җ�E#Q���d���1q�������PK�zMܺ  �	  PK  ў,J               179.vec���Oa����y�=^3{��e+[6�dS���M6�d�M6ԡǥ��}w�;���Ȋ�y
��<��T�"��������^��Ԡ��Ԣ6uRu}��^�4��iBS��5�k��ҒV��miG{��#��L�ҍ���o=�z��C_�џdP����CF��HF1�1�e��D&1�)Leә�Lf1�s�\�1�,d�Y�e�T.c9+X�*V���Y�:��ld���V����d���^���y����9�Q�q�y'�)Ns�m8+ϥB���hsI^�
W���T��&����r��<�y(�'<�ϝ�B��y%_�&�o�;��|��)�S|-��M�ΏB?ݩ_���PK�U��e  �  PK  ў,J               180.i��UT�M����A���}�w�� �@�����	$��A'�a6�^[n��9����V�~ޖ�/�7�׊�
� "  � �� h((�(�h�����h�X��^a����P��))H�ɩ�8�h�h�ə�ٸ��������B<b�|<�%A@GG�|�I��E�CMN����� .�$�B�q@��~ ��Nd��i��2D2
*:ƫ���� "��BFFBz����$\d<jn)|sT(O`|>�t�BͩS:^� t�7�$���L�,|��B�"2o����+(ji����ZZY��~��w��������5$4,<"2!1)9%5-=�������������������g_�������ٹ��ť��-������������������\ ���#�"	�?.D��p����Q�4P͡�4<�h����?�iy5O	-\�0���6���C��d���������˵`�^6�@�S�Ӣ�H`r*����k�%�U8���[��u�/C��X�~��]�g��#���\=���o����ƶ�ɪ����H�鴥f�ȒV������!�c�ϐ܃�<8�e 	�g+~Ͷ�vځ�^c�Lg�ˉ�G8��V��g�a�J�^� 0z�Z� 2�1����k�p�"�x�ꐫ��Z�P��*��{��\���;oU<�vbԌ�]9Lћ��:�͸Ҩ�]�c|E�8_�}�<
Xiǹ	�=՞qy������8��w�>����j�]�z��@#��[hVλ��q�o��=>M����|M�J}⑉|h��-���qZ|��HY���s�s��y�s��������1ɓ�6#+���IV��ެ��%z�^�ށ�!ty�	�1��W��`�R�T��@7���F���˽1m'�kU�A�t�4�7�4tcQe�.�$�����[y�j��P�Hb����օ;�y����gl���?C��H���A�B�~m���n���٪z<���R9�廞D�Ӫ̯+Դ��u)E��y��j�`��mgV�QѢ/�O���+!��B�����G��L%ч���(�^�>yy������x������;�U�ː�5��	�]kU}➘�p ��l����[|�-��<��a�cѓ}���7�Y�u=Jr��v�{1�������(���6o�k�<Y��{�{*	�e,ۭ�	7�}����HVs��E� :� W���V���=P9Q�t��&X^,�S^f�%��z�K�dZo�V�jg���{Io��_n%,:O��Ŗ��3�C�����%cp��#w2�VW�ȰEH	��~wM<x��\�/U6DjML����".V/w�f$�.���(��_���~5HXi��j'����i��<R�L)�ov�/3� �5\�ɪM{�14T��L�Zۉ�`�v�r�Tc���������E��u¸����a:�z��zN�P������������Y>K�쳤F�-ys�71�S�(k���W�:�?�>fT�F#p	�����s��;���/n���P��km	��F%*ΐ�'{f��ns}�t�y� �������+�w��*�4����S�	�5�6�x��=O�r����س
�v:+���n
�v��#
�7��:|X����q����҉9y�:�d����Z�G���<�)E�p���H��O�7�=7p��`J���Ӊ��"):o�I�=�nM�ǝU�H�AX��D�z�+�QF�G��6!fl���'��te����Z�v;��E��gw��i����F�	�I��IC%Z��~LGu9�ӹ�C����@ZZNR2�t/�B��0��1xX|\ʙ�hj$o�G��l��rC%)�D�?�P�?��!��?A��b17��r�!�nl֊�z�݀�Zl_���ö��|#9��A�'\Fw׽P����/~����nM�g$�S��}k���&�}A|8Ш�3���T��뉇R��2�gGzىv�U�<3XI����C�o����jߙo^��?�l2�:�3�ݙ�iz���Ӛ��i(�B@�@���_ig�ؖ[ u3��(	+@�>Al̘ߊ٥s)
w[
�T_f����/JEG�Cwk�8�o�>��B�_>iZ�H�J�u��UJ�3��5�n*d����01k�m(���?:�QR�Sa�0B�ƞUG���C;����_w)Q����m`S�̇Q��O�0�;�FqTI3S����u&0�_.�&�N�-��4����'{T6��kC�Y��n���e���qpc|��5zD��i'�)��VE��(���o�UB'�YϾ���e	��6������.uE��n.ǔ=�����c�x8��]�^�
�ci����gAiL��2f�#�6!�<���srR��sJ+�;�k����؎ި�������He7����ɿ~�)Q�XV=���4��(Z�X_���Y:��ꗿG*fU�'h ���-��3d9�����h�%�ڜ)�h{b���vo���b�9�H ��\o�~��U
c�4�Q|K��?� P��.���͗%x�&Fm����8��	���U��Gk�Ar�p(��k�����y� ��ǅ0ƩH��I�_��;�V>�8��ƔRNSͿw{��";�'(IF�F�>64�,�8� ��I�<�A
�/y�!�)����������Si�2_
��%Y�S.*#�����;�Y��N���ɷ�s��7�ORUwp�F.�»�v�oj��&2*\n7+���J������+���G��i��X����^j�-o1��&��䞕��ٟ|�UU(��~ܵ���;��5f�;D�>~�N4�U�Ĉ�v��y�hnҾ��6ԎN)ݩr�d�iP�&���(�Fblc�ds3��-3i���j{�oNV�&Fy��.�������|{��Z���Pk�^
at�����쳉}H��S/�ZHP���9J��GU��˲���3�>,튧����2:�t��Q�h/��3x�\"%�q�bJ�����"��I1ж��_�$���'��➉�;��J͸7�(9�&)���,�ufB�^צּ���$0�9ǲE�W^L&֧�%�,<�e�dM��ձ�~vEM�Su�1v���x�_*��h�:ɝ/��%mֳ�<��Z� M3��M��C��5�\*Sd��i�[~���3�֍$����d)�G^�>���h�0����h����ql�O�&���t�!���BR��糒)���1|]��q��K�D��H.���K2F���B{L��}�����������U7��]av�kM:*<ڋq&݌��E3nj�ς��9���;rp� �t����8)+�.��D�)���Rq'�d)*9iϻ�����T�Aw��g�B	�j��qFz�'�����m�9k� da�@DF
DI�k>��=S��JOlfX��d�
U�!��|�y�Y�v�7!��b�S��gh'���3�Hw`kC����)n�,��F����.Ͼp^C�6eφ�0�ʛ|�vhO�Zb�q^([��]��2���O9~@��C��ɑ�?�0��*z�	"jzw�☯�p��9�4b��1F6��^O+t�b�:>
p�*����Z�Y#����9
���-���r��E�q��Kwݝ��^�+�|:Ly�������δ�.���aw���r�Ljɘ��Q�ZLL:�i���
p�;z����bi��~���-�(N�0����r�G��W�?]��(�ie)5��1���8�$� {�����.K�G��k��)8p�SPB�r�	)!��S��B�T���JøKNS�������S�� K��X�M�HA������d�����h��A�@�J^7qy�O�O�5�{2�\�=Xg@�6����}��o�	�Q:�2~�a�l五w��<��VN� �6L��'ш�3����.k��Df�[�����N���r�3�����$%�	��5�	�M�����_پ��-ۗ"��z�\ke"��~ɥP���絣��}�zsK}Ҝ$��s+�Ж	U�C��<��R��B�Y���9�6�V?�~HU�����o��x�#�����s�)�,��Z�d���,t���������%��U���Y�9��ݪ�'6S�����9�)GE�m���銕w�BwzՊ��W|�+o#��5n�a�T�8��`+��&#Z�u�(�N̵�$ڲ�ܚZ64�m�M�����:�����
~�;]4k��ĥ!��/��Y�0��*j$[�nj.{�p�K�k$�;��bX���!y��V�����~��P(�����@c٥����@w '�G��A�7��������܀�b�"+^K���<o�O���*�~;N����\y%.8��.c&?SζV����tp�N[�+w�!<	��G��j������%n��˛��!�El&8��
V�q�mF�S"�B�q��[����Z�Z+&���������џ�
��=,�G�HA���|w�#�g����E��gS��A�����08@A�i��a�V#l|'u���G'�]��U@d��ݖ�5�[��ĘY���L��<;Y+.� g��s��&R[*[ڻyCf�q}���X��,'����C�25�.�L�SH�_ҼhFI�K��|�ʯ`����i:ޝ�*��~7�B���gG(���g$�諝O���κ���q˺h��ݰ'�tCDA�{���B��lhm�	l�ɸ���{�t/7���Fh��fc��U��c�8�/�W뚑��<9h1S��E��Q�b������m�$��5=�-��jM����`����!�����)�D~�ާ�{�o�Ƅ��Ǯc(��j��J}cNn����x���Ԏ��u��4Ŕ[�2إ���^�o�����w<��7s�f~Qf���>�����Ո�	�O|f�v�7�!��#(����]W��Z�`�"0W��M̽�T��7��x7�ېʿ���VI3h�.��ɃY�����z7P<|���H�u��,�%�p5�]/=�׿x�����,�SY@^��g]����δ�pO��N�!��8i^�/���~1��Ir[ܻ��O��T����m�֛����I˴�J��nq��K0<��8s@2O�9����E��i��'w�MC��X�1�l��~&T<����"�NL&���F����]����eH�@��8*(wOO��Rii#Z��b}��
�сN��B�$�ٓ�Է��#2�bZ&���N�,��!�0�=�$x��z)�����%�]!y?�\��VD�&*-�	vS`��T����J<У	2�_ϫ�>�k���V�.�J.ns\||4��)h�X"h`��e}���� ���]�Vp��0�������L�����H������*=G�U�P0���,����"�Կ�6bL�D��
Ա?���.�ՙ��^Rg>35&�uqy���w�QwHr��k��-9�<K��#���Κ��$��e��|�Әvj��:�q�ky/����4�;�����{���ʴ9b
Y���?wZ+��9;
�_���mu|��m(�Cؠ��U���W���
����"S��\�$��ڑ�t�o�m�'���j�d��ޱ�й��9��9��[�^O�&��&	�[f^I}(�}���α@�y)��1
��Ϛ	����@"���a*z�+��D���v���nU(���1��� :�챢�*'����m�����B(';��e3����5mB�� e5g9a\u��ü������`���\{d�b\��q�-vE2xd�}��^�L�e��^��E�i����ٔ~�)E�qV����(�(�G��>3�/R��n��US��(���ᜒ�.9w�z��<���O�O��Nƹ��h�Ŵ��"��?�ݟ�*ѵ�7���@�@P���v�vZ]�Q�AI���ƘK�1tXU�^D�7�s3�%*�jt��*Wc�;��ARI�L8a�=V�S�sU����X흖_�����ډ2���!�Ě��m�ζz�����F~�`���+��h"��dʳ��Z9P)��^� �8y��*G��&�񉣂��9 Vq����3���=�x��1�$�{�<Y��IT�n�{_�Դd���s���=�ʸ�8�%���������n�ۓ����ڻ�Au�!4$V&������1�=�p@q��c���+l)a�|�=xQ>�Qo0�S�al��ĚS�b&��<���fe6��@�b=��L�btp�3r�&���;0�1 ;�Y���U ;��8��/�pK+��@Ƽ{��kyo2w��tCRUq����Kz�� 8���#i�YҶ�i�]�3MȒl��&6j�p�����i��&/?�?!�U)t3U��vy��*!(w��d� �v*���-�>3#�<���=l�f7�h��(,��[�>���r�@!�"�W��!d����mKa��ҚYG�����%쑕�(�-G�,r.���E|��VW����)Q� �9�9 �z�_���CM��V��oI���x#�]A&�����zT����ハ_�`�
X5����F�R���l3)����K
����zy^a�r�ha�3��b�F��X.T~����$��@W����e�H�J@���N�ڽ����ŝֿ�g�/�.^�ZuɅ���$�1���lL� s_Y�t�$�	b1�<���S�]��$q��/tq<F�r_�9I�¨�_������.ux^�3�_:�~�g�%$S�-و�GG2��ܶh����r\TN���Q25!�xPW���=k������D��;�ٜ�79�!�~�6���a�2�˝e�}�컐��#�q�&8`:]�e�[��yX� E�L����X�Cb{�&K�$v>C�Q����_f9+E��r��^��{��X�"�WdOg|�:=bD^��0���{;A�^+��(_ڭ,�H/���-��Ua���\�n+o�S�~�k+�q�����b-�b")*�1��%�{Ǌ�M���R2�X�h�����0��`G�X<){z���B��z�i��j�K�Rz�&"gB5�*DF��xW��c�%�.z�Z�JyZ��6�Ҝ���b'JkO����^�]�'{�PsL5��_���n`{�	�	}b��]��X����^�*����],�)���+E觚ڲ���^Q~�������xk��">D����w�] ��s�yu�yVDн�^N*΂��q��[�����H<����iL�O9h�f�/rr�|�+0� �-��!|vo���r4BO��F�?�.��Dt���L��#�4��9A�z�[�b���V�����NDɤϔ$��mn�@Vi�e>p���t3��Yҵ~߉q�nτXt�-m��o��ޞ�r�|�8��E� �����`��͒Z}%� ��c�Z
��Z5Xm���'�7�5g���/9Q8np�$M����cH�ntE�K����'�o��f��Zb��;�
t��՘T��i�T���c&��:��L��R�e��u�$ �xۺ���!��{�9w�%-��cş01��e"8��ʆ-��:s�d������XD3�M91��&Ύ��>V� ��k{��(Tży�Z�~��6����a���y����>C&p�O��� �	(唹,�Ir�ג��B���i� ���ᩫ��������pvwN�ձr�]_SҸ*O ���}B���Ax,��ZWer�v�ܴlL)q䟫89Sc�:���G92ƿ��l�)<��2��u-�Y�:g� �̾w��eQ1���\A�c��Pd	q�N�����8�:�,:�`M�j�I�/m<�g���t��q{����9�8����8����	�P�+��i�5��eFT��lDG���{��{f��T���㗔�#���%�b˷��Ud��i���ܘL��6���J�G-��:�}dQ�Qk��� %/�p�R-@�M�=w����н_ʍ��m�\�Yh:7�!0W2����<�ĺႢ6SzU�[{&_��o,�>�/7�%���	Ҏ�/��/�PK�d�F�  d   PK  ў,J               181.p͔YT�W��/#�fb�U�A�!`Тm�j
ȯ��@�HS "�@5�(�P�08�)(��2E�BTX�4��ᦕ�]}��W�Yg�������|���@ ��~|��� �H��%�b1��`F��&ϵ����8.t�8�PmmiK绸�1�L���r�'33��(
��Z��Z2�m����	���� Bq�A��>����S 
�#�&(4Ƹ��# B�����$c���x{7���Cd�)4���ZOZ߮q\,�MA��-,����9��/`�/Y�������X�	ް�3ަ�͟�G�عkw��/��<��Դ��_�����8y�t�������%��_����z�������Ʀ���;>z�D�z�����`P�r��ظvB����ɩ.�������� 0���!�3p0����En�!80�W�^�GQ�א��hsG�����d,�/����\� 
Ã� �i�I���\��,��"��g�VUt�ʱ?d��Fp�Ń{�#��N�_J�������xn��H�������J���Q�����v6i%�&M�;����ϳR9���*�X#���u[�O�$��JW���,�Ī��wr��r�%6�	2�� H���8��R&tU<�l�{R{#�	��虽�L� �<Ƃ�ϥX��CA.<�M�&r���)NBI�����wk ~���o�t2uؕlS�`�"qұ��� �0�K�Y��0��u�%c�U�]GdBX`�>е���[�����1���ռ�+wv�6ʯ���u����c��Y���|�E��)�B��c=�mN�R}N�M)#zo������I_��M8�sRI�Ea��<J��E|�T� }����ϫ�+x�WZO��7�р,H%�ʭ��8Vs�Z�fWd��]�f�X�kE�����IE�YC'[��F�g���H��	�c?}#~R��Z٪��M[�ܟ���B.���C��1��,MY��|�r�5��/޼�����KV%�X���I͑E�*��ୄ��A�7�R����FW���e]�Ϙ��Ѳ�,\�s��5�[����ko��y��E*����1����;{�ir-��%�2J/�A&r�+6]����-
u�r��5N�]{�n�u� ��y�T�h��Lއƾ�mQ�t@"��t2EM].T�2}.=�+l�S�Q��kN��,�y��be;r��:!#�R�r:��Qq �n�u���D>M���^d��b���YSy'�츰�4N�}(
��W�FEO�q(��Q��d,�حΩT�B��n��o��h�wF�Tj:���rOl\��8k}�$i-Uw��S�h�����	�Më���-[��s���Re�7Ò��R�S�M4��ƿ.3 q��O:�Չ�%&}�ԦGJx�Ŧm^�����UՄM��{��6s�lM�����@F�3NU>+>����#��r61xV�3Q�|�E�;7~k����:�n��n`�2xgq�e���[��_-J�O9=.�J�3��,�Xf�^صy���y[GG�`�6xQƩ��f�Ş�/��q<�!K^��s���*:� $��/�+�6����/�.�4I������5�D�è���}Znh^��[���U1�w�UT�.��Οo����e3RD�s�����WPKdu��  m	  PK  ў,J               181.vec��a��3�{��n�^�c��Vl�Vl�[P��Vl�VԵ���v�G����p�7"I����y
T�
U��%Q=)DsMjQ�:ԥ�i����^#sc�Дf4�-i�}��1����@G:љ.v�j7�Ӄ�������*���~��` ���2̷�7�<�QN\���X�1�	Ld���T�1����3��l�0�y�gA������,a)�X�
V&�JW����c=�Ȧ�<6������`��ߥ�)a{��~p�C�HZG��9�INq�3i�z�s���\\��\�sU�q���VV��z����>x�#�y�Oy�s^�W�捝�����^���'>�%��Ww�-��^H���W.������o��PK�줔k  �  PK  ў,J               182.p͓gX�W��7o&!B$(`����	K�1,g����:
�(�*��1��Af��Apm�Y*�"�-$�Rh����B�}z���t�s�����3�3/ uw � �<�L��H$
�@�P(��J��b���5��:zKuu�D}�9U�ДD$�XƦt��G�YimionŰ���`0�XU-N�Ҁh`��c�.�G�N@60<���J@O�'���� 8�BcT�ʂ�� � B �pe��2��tg�7 eN��9��&�*����$'[F�bT-���1�Pi��+�,k[�j������'���y�}|��CBö�عo䁨���㎟�?y�4��0)9%��(M�+ɻ�_p�����w�*-��PYU]S[W�����I[{G�˞W�{����P�4<2������,@�o�\x%��Y.5[��#�ȅ�\T@���e���|N�=��S�Ѥ���xi��E�H���b���`pu��4�����&>� p���Z��d�
dиӧ}MDY��-��}?��M}�"ƨ2�+;�6�k����Ef�EԀG[��-�q;=��E����e�	\�_j��Md�[2�3$�v�H�� �o��Ӯ2<�v �A�)��2�qc]︸�GΊ���=��
��r�����҆'�)B��JY+e����!<�K��\z59��1�:��<��l�k��Y���B���7VQDJ�u�>ц�;;*��d��ës���Vby�{���LX#��	�6�%����l������z@�{�%�Rآu�1<�����m���ȰM�.��f4g�-5�+7p^ �C�K`�x7vp�o��bc�����}�C>#.0��T�1	�3�o��__�Nr	e�_��h�
M|l.�nP��c2!�x!��Z�]ʽc����|0vP��ŇV:��" l�gl2q���xښի�E�|Z�1��!(O!��zEC5� 	k6!K�LU�>ո]�RQ~�+�	�|��>X�;���D1����ݢkF�hc@1�6��3�=$�Cѓ�<��������D��H���[R
�Z�<��C�K����1�X@�R��^V���8�;�}_�p���T�)m�4\o,�fқ���}��!:��"Qe+۬��͸�O�P�I^��&�&�f���6�(֢N�ix����:T�����׿�j���\���s�])��W�|6�)�'�R5O�ʚ%э��g�
�U�\j�gdv�?=��* j_�=)�i8;��㝃g�]�E���m3G�j*�rnt�T0߂��,����&0u8�#u(�4��T]�q��� {�R&����]�$Wk8�3�4]�p�PE�:;�w��녗V:K��!�`l�F���x��'�n��=�"�wNߌ���[;U�EOo��c�a����͔/���� �k�֗��y������ʾu�B��n���[i|`���v��%��u��{t;"�i��d�c�o�ֆ��=�z>���y��v����*J�m�F��;*�N{e����@����'�j}0f��48s�f��"��޹&��ރH�l� �((���α��x��>��6�z��q�i�ם]���O+x�J�Ks���g�R�G
];\��J��m�IBSl�3�`U�eX�� `�@Z��������+9�:YDrt�O��*����E�:8��PK�q?C�  e	  PK  ў,J               182.vecчˍq���9Ǳ�ޛ��k�-�l�ɦle+�l��&�l����s�t���|�ө'"���'G�2(K9�S!eQ1+D%we�P�jT�5���Qۮ��.��O҈�4�v���iAKZњ6���M{�@G:љ.t��Si�����Eo�З~�g ��Av��CJ	��F2�ьa,��&2)��d��T�1��d��|�ѹ�c>X�"�$+�����`%�X�m�ѵ6�t=��&6���lc;;��.v��3��>�s�X��z���(�8�	ߟ�S��ߟ�s)����^�
W���T�z�[��w��}�<�G<�	Oy�s^��敾�M�o����G>�||N�K��k��"�w~������PK>�ٲi  �  PK  ў,J               183.p͔iT�W��/+IH0�I � B�"��A����H�U�lR�`A��`AFY�"�FY��i����	VYJ Ԓ4x�Ο)�̙�������>�}�U(^�lW �  ��bpT$��D"Q(�*�����hj��tI����d��	�h���>}��K+&�I2�s�e촰f2�Q(�*F���}
�?�w Nt��� ��P�� $�9��� ~��H�L��   
�A�pL9{J9�ppM��.��0�(�H�.Q1�]�H�ꚣZOA��7uti�M�f�m6�m�v8��\���ݽ�}��������а#G�c���şHH<{.�|?]p)'���y�W
D�o�,�UV^Q]s�����M�%�hnimk����{�?�|���蛱�ɩi�laq�����k^  ��SzA`0(��B��p08�
����<�e�HV���.�jD[{��w�����4��G�O,�2�C�^��*T���v�(��8�?�)b�B��0�
�{�C���(����5�j>��\�٘�zIOx�@I�/�J�ș�e��t,i�d����Fq�;kr�>�[���۞�7��<=�c��p��֬�֖�7$���4)T�Ћ!�v��W7����|>:�Uؽ1���3�E�C-��4�+�����r;-� 푋��T�0��Vv<���Yq6g��U�HJ��E]o��#��H$_�ǫOq�gf�]A5��a�tљ?�^]�����ʕs!џ���I�7�|�Y+ ��_GE��%D�O�������g���-],���փ�O���;���T��������=��8�V��������2חv�n� �n9]yu��v��j�o�Mgc\�,�O�rU2��i�4i�W63�N���4�������9�<9,<��o�5m�2sýs>?���������Ujɓ:N~��䄽ysW+�� ��</����Ԋg�+�Z���F��,�r���=
@=ˇ��D�_G����tu�d��Ggn��?������^c�.Ug�����-J����.�t���Z��.�G���}z&˒$T ����i����;t�O���7�p�����@�K"�%N<܆I6>.Y�'��-Y���TT���2�}= �Tr̃3�ô��� ��ƽ`�U�Pu���'}kh�%*��V({|3"s4 4 ��c:b�O3��װ��t�H �ｸ;[]��$��{@�ĝ�}��k�e�Ɋ�C1w*�%3by��5�"+ڀ%0g��.3��?����d�^_?X�i�̲���=G�W�)����?��NI����6�g�^�³;� R��V��~|��p\���4���]�����7>E���]�x�o���X_�;�h|f�쥿w ���^�?��84<Mt�>��U��7��nj,#L��M~�»�\x����l����<� �|�[�{����Q)A~!���r���$E��1�	;R
���_�w6^L�]64o��!�����\JOk�	Ls7z�q�����1�Y�X<r[]�(����fD��~��<'��5�y�zϠMo6g�4� M�=(��C��Y��s.��א�͛�H���F�DQ�U�b=�C�-XM*�����~2q���ι���+A�SI?}K��4v]�xB�Q�����1����\Msګb�	]������-��/9,�F۪+��
PK!;�`�  �	  PK  ў,J               183.vec��ˍq����p��&{�e�&�l�)[��&�l��&�?�>O_�NW�O缻;?�Y!2��Q���T�"�����bW�]��Ԡ&��M�<���w7�!�hL�Ҍ��®���iC[�ўt�餝�BW�ѝ�qO핊�ۮ��/��� 2������J�(F3���c<��$&3%+��:���`&��������,`!�X���,+�r]�JV��5�e볲ؠ��f���mlg;��n���}�� 9��qX�p�c�'9���z����<R!.�%.�W��unp����w��}�G6��	Oy�s^�W��y�oyW��{��G>�/ޛ��,�R|/��#R��W��w��oJ� PKH�yd  �  PK  ў,J               184.p͔{<��ǟ�g��4�0LSL��6��!�h��Z��d���%4D��uK��$L��)1#�:�k����ے�V��\�9�{^������~���y���H�$��F[{[  �t�Q�@!H�D"�h�'���Ũ*(��x�f^]}�P{�����:�LG;��ؘ�m�ku���1u�!4��Ũ�ɩP��o���<�(�p�h P,�B$� Q��\�?
ap�����m���@8���H����b�PdCj�p�8�u��;����fIFާ��2��UT�۴��:��&�f;�-l��m���;f��~}����@��gBφ�GDF%$^LJN�ľ�������_Pz�������f}C#���m��;���']��������p���kћ�S�s���}��� !���腕zAa0�\��@�W`a���5y���A�C��p��y��4r�U�>�'��d,�6����쏉��Wf�����!��X��v�K��q��G�
�?x�=}��b``�so��T{�-�2zhKIX���nk�,�<�v�č�+`�+ tܡ��wͪW#��t(zqb�� %?cr$�?���6�k�C�o�� 1��W�M�v�C������Ŵ8oۧ�\�Zbȅ#����'~Kq���-�+��h�(��7�BX�R��Tm�Nr�!]w	/Hge�ˌs��~-zc.jQ���η��Q�X��w�gN�F-�Sa���I62�8�@g�����\��m�ݨ���O�j��Zy/fF��]-m�E�E��G��yN>z@�u���`��7dȄ��Jq�R�Cp��
���&�1�3�+����j͵��u�l��P�Ĕ6���y?gX�	z*�o(�}+P+g;��:_�G�F&D�<�'E�����?J�W�kx����J��^6�v�/�n9���7�sp)(��wэĶ��z����i������5�X~�����ZYo�v�R6Y��OE7+�zc��0�P|���~��pm:wֶ��Q�𶮼��+66HI����2~�JP���>�/�l��p���Ch���$�e?���$C}����)ؖ��(��?eM=)?�̓v��cЁ/q2�b�r�"�=vH	�5�[�+��?��J�g���T�čԑ��q��U⾚��$�"����/�m�{�,~�?xC!��7����:��������Cޮnc��&_�~٨�=�G{��=�{�>��#�����g$@����h9�t�G�����a&r��[�������1����c�7���%u3tP�\za-,�R�㏟�5��æ�z% ��j��<Wq�h��6}�;5���ٙ�z2�qs���ϰM��foi�k�yk ���d����K�ʻt���.���ӝ"_���}c�{�e���)��쬴K�����H����QI)oG4,�,��ԭwMK�o�s�¬�28�U�]E�^j�p�y1 �� ��a��R��3��˙ӮC?�����Y`�=:�at��s R��Rr�׵^�,��CS��X��]B_8�\bR;f��۫��f%���I	�}Tei�ܨ������ݤyb4�%���J"�*a@7���}���S����P�a�����f/�ekT�G+�`�ݸ��`F�!H��<i|�3iF�����=}���%̈�O�J+'���Y1BG�h�-�̇���X�,ߕ�e�p������'�J�d��PK��m�  �	  PK  ў,J               184.vec���Nq���y���&{�lʖM6�dS���M6�d�M6�yn_�NW�O�y�v������2�u����@ŔE%���*T�թAMjQ;�QǮ���i@Cј&4M%�̮��-iEk�Жv����Dg�Еnt�G*��v�ܽ�C_�џd��`�P�1��d��X�1�	Ld�����S��tf0�Y�f��\��|��E,f	K��X��Y�JV��5�e]V�����lb3[��6�����b7{��>�s��y��0G8�?>��9�I�O�i�p�s�O����T��^�*׸���z����.����<��<�)�x�^��浾�m��;}�>�Ͼ�/�_)���)~�3��|{��R�PK�3�c  �  PK  ў,J               185.i��g<���w�^"Z,�%���%����$J���UB���]��B�袳����-�>���7�Žw��9�s�{��f?�_��T�P 	  ���1  )11	1)			)9%=%%-5=+3���a��a�/�@x��ED%$$�<�r2b���%��s������LE�p��?�@C
T䀀�4@����I�o����IH��)n7�� A B!�7�� �!��U"�ӷ&��N/�K
S��ɀ���)n�BF~���������/!)%-#�P剪�:\C�������������+G'O/o���|�B?�����JH���������_��ZXT\򽺦������������W_���������������v�upxt|rz����?\@ �?���Es�E@H"$����6�q��*�X���&�W�ϭ�IG�3�x�&��)��u���&����"�_`��k@	�&DP ��D�����$$�H�;���q
N�w�nV&kI$(K�v�����E�QO���Y��7���W�cx@ �� �˒��Z7�����w�&�R�k9��`�%� o��HV-�b�Ь�jOy�Ri9~V|�p��~���m����s�t�3o����ʕ�Mw�R�P�N�Qo�&�e~
OvC��T��}Ɏuj�J ��'��/Y!͏��ڬ��y��|�@�1�&�NuK㋝~�j}x�cݪ٤�PU|�����R�rl�NF�a���u'N�h<�1z�v�_�`�m��)$��˲f��v��r;6�����>^��D�Trv��b��Y訸��s]R�:N3it�y����~���ͫc*/�g�ܑ/��u����+W���*�����˺+?wm�%�m���tn�C��L$>�}�oߡJ�ԭ������7�_�j�rAqL��r�j��#�ʫ�v0�V��\4�d�ɦ42ꦠ���#�>�ZfRx���Ή�V,&��zWi#��)����ۃ�r���X�2���c Ɍ����^�9��m�X3S�����$�~�G�=�-S���L���+=OA3R M�D��.j}�}�n�*�J��@&�^O�xi�uN}��?�F�>�W ��#��r��S1�/-Q;$B'�����Z�c�U�°���#ۦm�>;��i�Cx ���P ��3+����M�}��=9ͤ�Xd��S8x�0!Ǘ���,���ZHG-�b��R��^�g[�8��s�w��ޏ{�D�#��.�����;ͼO�O�ۃ��:��e�,�(���'b�{̹��V�|η���O���6¤}�9b��D[73Ƨf&x8����k������tq��͐��1<ߚ?���X��*��ϖ�i�
,'����L��c�]����}=\aC<�WM��B��@Ėu����J=;���98�珷�
�H�=2>�H35�KR�s���9��󢯁�N�����?e[�)Fկ���w0+�V7����KF���	�5G�Pפ�WNr�Γ��I9��|���&��p2u�v�T"d:����Vj�ҍ�}�ljǝ9뒬v/�a֊�#:��I��`(�w�@Ass��R=��2#������i��c9Y^�70<��b�/vAU(tXX�g��/SzI�
��;7ڵ[�Ә�	��2����<Ӊ����9��(��}����=��� �,�|�NEPB�AV>�R�W�
.�|�Y�~w��n���=�����8?�A1��NSܫ�5Bbug�w"��yÓ$՞\Q��2��ue;Ys�oyQ*�l,�r)L5_
��r�&��{�����;��uj�g�`��;�u���Gg�����n��Aob�aUx��q�Pes,�$� �=�*�v�8a�<�[G])�mԿ�Q�Fx�;�z��W
T�u1߽bB���z_���O_�Ò4� ��<��aw�C��ւ�c0��;j$L��'���W�c�/s�uY@�>��l���)h�#kk
�v���Ul��2�G_��a��9+U��j_�u�'-�y��t#I7��_��3ع�����,{���һ�^g�FEF�x�x*��P�GphyV�&)�L������=*��b,0N�Б�%��� A�����:޴���Z�݂2צ�1�`��� �����T�J�@�³�O�DD�F5���cZl�H�7�����"H]��)�������@��� L,_
��{�dZ#آ1z���Z�sFc?ti�s�����z���#����:Fcǭ���.ۡN��Ƿ�:ì�J�f��ۓ�;u+4�%�3ސk��)Ml�:|�$'��R�����`�ć�>��1S�h��H.���Nv�?�L���g��
�	�#�o�d@�r��Q�o$�Y�������}��ҏ�~�D����j�( �lRi7�̣�ݟ 5ۣ{�
ڱ�w�L��ْl0{{Wt4^zÞ�lM�ɍ�����bʅ�j����k��e���J�;�Q2z�-:�n#�z��������I���y����n�`?�@��,.�\J�� ���N�G-y�����S��KI������,�����B*&�SU/s��������^���	��$��4Y����4�铝�n�7�����w8/�������,-�}b΍�Y�О9��j���s��+�V��l��F�Â =p�;�*&X;"}N\���(5���_�<����̶QC�x�u�5����ACp��2Q�T-7B� l�c�ձ����+o�wE����+,e7�za���y.E ����x@����0�z�A)�
�d0M�ˊ�lK"�M��PL�N-a�:�y�(߇���?�&�o�9�u����4��¾�K�����h���|��!�_Pc�����@x@,����1�;G��<mʪf�E�Ƅ߼�=KY�Eu��!�Sv3�	;7j���ύ�Y���5�dރUaء�7FR)����Y�x*�Eo/
h��pB��H�q�d:#��T�[\A$�Y;OlύH�_��|5(es�;�t*
ɰ����5��37�^�F�+�%��v��k��V���Q����)̕`��G�ß�"՝!?,D~B�<��D������l.��,Ȼ�t�<�h��ct����@]MQ� ��� U�̭	�O��?�,�q�6��|���_�Z(��=���L\/q����r�ā��apcӤ��5/�e�K�Q�8��إ���ѭ�9X����H�� �s�j�1�諊�r Z��,��r��,�ک�ɇW��0̛bZQvSÀ�u�� � [}�\���_b�,��^N=�����%���R�}��뀧�OKc��-8}�-pk�fPM��
��:]���$Ɵ�)j\�Gއ��m�&[־�Vq��9�)��'�j��H� %h�z�4�\�$�?e�OE��~�I���2ǒ�'Rq��Zz��Sх�����՞=�;i]�k��l�� ����m��slފI���Nܻj2�xP���3���ej��׎�Թ_LSbi���û���[9�M�������>c�>�Fm~<�)c���kW<�^x���O|o4E��j�y�|��'����I���,i�@�?򐅖���+x��+���ZD���7F/O��X&��J:��dY��NV��P�	�j��|��=���ߨ��t�+�r�{���BE��d�rO�&�ۨ��ޙ��
���$}[�w
�;���̍����š�C�M$�bߔ⻽q4s�8\d�a��K�����C�M�7��y���r<r�`.F�gACU8���k��w����d�_2U(N�����"؄F�q�.�E���WwSi�i��_��딗^�j��uI~*���9Ah"%M���v\B��b�q���mF�R��	�➱6W�z�_Ë́���BǣR����@����d������N��qB_�lٿ�^S�r�J��j@��s�q��lo��d��:�K�*�u����/>�)k~21RL�>�o�Ɨ��g@�v��#I3�.�jv���6n�"�h�1����6����rT��4`��
v��(djh�t���Ծ��A�e���S8��S��y��~L75F�Vn'pL��ت��m�I_� �vG��ָ�������o�qqE��Ug��~�8��'������pZ�N �!t[���K�j�4{�Z&�6b�ST���[�X?#��?����]!�uEX5�#U�=��B������Or:�c@�ӒT9ܻ�;ԩ�W���.^��PKx~�v'.��/��yl��N&U���+��3E�����)�,P	�=?��J��O�l,`�{�'�:I�[Z�䋍.�P�]�mSw����Pi������BZI�=�k(,��<}�_�����H�T~<@�B����S���pn>�+��K�`�g]c���mB�/V?1�	��	S�K�JO�8��k��@5��,���ܭ�˂#?9���zף�)��N���. t�ȇ-�M7�����I�%��w��D���A�q�KE����HKhG���%Q���U^V���-V�)[�<�(��QQ��8��$���7�>�7C�k#;�alF����r<�ƣ�u��%���$�Na�_��h��q'�G�_���<X���p��t��)=_��v���G�sz���U���4��� H��;2����������c���\��T\UfA��D'V
����Bݍ?�Ed���X_EZ5�/�V�U1�ml�(����bX��+:��3�pZ'�򇽱H�ܩW�R�%|^�@8([$L�fQ���j�zߴ:�6���d ?W�R�3���H���>��d�(D�H^�4�w��s�ϛ9��_��rc�:A!,A�Ӡ���yl�>₎�� L��ל_����&�M�Ҥ�w��/�ł �-��}=�J%3o.�f��;?�J�#����h&��9@��z�t`4�7Y$������_�� ��	�HP�Lߞ K�s�<7o���z!:n�c�gy�����K�5��IwL��9�b;������Mʽ�ÉK�2�Ğ)v͏�_��ر9W�=X�񐃛�Ud{��y�ғ{�NQ*��F"D�V	P�(?CM�]4�gjU���6����ˬ�5��f����c���(���D��c����h�sΈ��?m�>�1������>�������^��n�IӜ?�����t�\����6|�-�k�T[ ���8����u�z�?0�b�SCr#� *.z��J%�����ԉ�+�A�ʲ��֏�l���t�p�����.v{_���3\Ic�s�_�H�]���6ewG���A1���h�#�^G	(��P �9O*p,����t�`�ỳ�������sV38%}K�|N��R��.��I�x@�u% ��p*`�#��H��-��N�~���]�����-�א��P��Ps��?	W�k���A&��];���HͭUu�2����#���[N��X�BL�h�=ͮ�Q�8G[�q�3��v������i�6�������Nv�X��쑣

�x��+{��+N��t�3����6�7��g����t*g���)�Y��I ���-���7�z�b	񛘛{��2L/N�&�������_D��I�/�,7�=��yˉOi)��G�ۆ�'z�y!�W�����9q�r����)~�7�cx��ؙ��z�����'�2�8�#�ur.i7�m�Nu
���'�t���A^����L��g(�����?�h������|�*"P9*?����7��Ȧ�o�`\"S�#��,m'V�32g��E��u9ƪS�O3dYȳ��pռ8��ΣɦBۋ�t���>}z��^���vf��YԿ�<�іk����S��������0�j�@c|[�_6�Ϭe&87E��kNb�<֪_�}�,6�c�%�cvM��ެb�}#�[�;�oD4d�%S i�a����w]/�9؜���+U�}���B��y����R=�[a�Q���U^/� �-���\������=�Ŷ��CKÜsي���*J�_`;Z$����Ր�����S�� �Wqx�c<qt�߽�L��@'r��m��/(����#m{�*�\�h��U�\%�G����{��p^\�v�pk�h �v�މ)�(<�C���g����Jͦ��s��ݰNה��;[����ܵ�)G���${�X<�M2~��yvֽ:��O�Ul+�ڻ�Pr6��~ş��f�.�
���˖����Xx*Ivlq&��&*�C��YC'��]aM#���Q�����FD�Φ�D�拢5+�ҵ�M-�]�"�V�SlH��*=%_���F9���P?�e�=n��\e	��F7.\V�и��)��w{���47Ut�;�j%�u�݈��Y��˺߷x�$#������XrJWv��� Ι�K�X|*Ŀx�O�K!Mw�Ȏ���ά���d��u�)�yA����nv?�Kj�=�"�P�,�LK�̮�V[�*{8q��E�(��ʁ�4hq&��,���V�x��@h�^���o�Q��p��=����Й� ��������"T}�u�M�KX��S���%;�}z��V�p)�$�G�H��w��_)<���k�h�xs>���cA܍6����9��
hRi�"��q[C�c��Ò��0A�����5���c���͕���Is4��=�o]LҊ̔k��q<*^�$_e%�^�'5,���u������>�O6��ϻZ fNa
S�PN��^T;t��)zԓ���Aͯ~�wsȢ�E�p�o�G�~�OV@�0>g����Th�J�t�5yl���L�n�cB<r��b����ʛ�8�H��b�7z�VC����s7�2�$S�\�`:���顆L*�E�(Uxy0�&}���Q8�MM��9�Gܪ.�����dV�wt2�Aq�nȇ������0�&�I��*^0��"���
����P��b�"�����p��Z���.��WN\2
�pC_`s��!��)��?�΅�t5��9�|P�e�7��9��I�Ƣ>�Mako��;�6����뢖��{\��~J�Q�k~��=�@�q���̅�@���������p�_�J<�|v�և�`���	����E>6�����0����=�'�`u��m��Զ�͈;5m�Hs�mx����������ifwx�_i٫Ȋ&�讒�8�3ي��
Ĵ�g��a�`R5��-�{���cj�ށ/z!79r���t �6Kr3 %�)���螮�,7|,����{mj���d����%����[p��#o^jHf+�X����5_��l�c>��vRA�C��g�C����9�"U1���.�T�c_f(!���=t8����0ۈ���wZ���v$��ci���������%Ǧjz�����l<�Ȇ�	9�v����ѝ�=<#[5\��QKQ��^�I8����n��\V�u���:>_���e�l�J�7U�Muճ��Bѯ6�fk�� ��J
E��6B���Q aU�MG��qߋ�̳'�%��c*��6�E:��!��6��Ѡʹo�ߢ}{�0��*��N��A���z;䆩C����*����>��o�*3�V\�l��7��1�E�5_~�/8:@G,���w��B��}2��b۳�kqӭ@���7����"��߯>�M���=�VCW?α��%�tH�w�w��*'���g���T>��os��6�n�7f]Q�U�ݛ?��ĥ��s��}�'�7]�[���־ǒ0�ٛ��M�m�ί�S�6*�،\:!��6�q��]N�[��I��"��{����s�/!������EA��˃k����ϗ.�%;gF�
Yj��:,���$.zx���Z������c���T����͋�/��TU�e��I�:��E'�~��\+X"����C�m��^�Nf���'�}W~������PK�Wm  �  PK  ў,J               186.p͔{<������b���a83�T��P��-T���A"��ȭC�R�M���0��F:�����E��h��dԺL��2sƾv��sb������>=���>���}��>�K`�vGG �  �\�b `*WA"�(��*��VSC�jaV`�HD=�l��J6ZM!hLW�cXZZ��V�7�oZcai��D�Ph54^]onH04�Ӧ�h��[�(h@4A�&�hH�:��/�j 
�#�*(U5e@�J B�������iµ��i�5O��P�V7j�~:clq���R���u�L�B����\�Ն�V��m�N�.�=������k��ÁA�G�r��G���ş:�r��T^F�Ŭ�An��jQ��e7�q������vSsKkۃ�������L���xdt쟯�%��oe�����8��P�7��\�J.�!�@H�b�&n�@hٳ�~�#�$�V~au#�b�{F�穪��尉t��?��_���o�~ ���쀙�4���X֖�GaL��9M��M�k��
u�j�8��A$�AN�f�X�\s"�l`n$�Ӟ�S�u!� �� �/�f�p�:��$����Cr(H�]���[.�hd(��x0���IU�T��I9�e�r�����7��E~{
���z���z��Y���Kb]Ľ�@t��$|A�R�t��ĕ�u��h��d� �i�;��̽��]��Q�H��n��H�1��[g�;/LZQ�}�rH��ݝ���ߋ�Y�FK��m�h�0!o8,�v1��{^N��7�V�cp�����[���G�h��!�$�]��g8�z�S��!)�g�+c��w���]$�xb�<�>u����-^^}�G+�R��S��U#9�4�����"��2n��gyw [��9n�����w��*W���6S�&��R���L�t����_�<�5?�9$c�V'�#�ۗ�^7L�~1 (
9x�]�8 �����Gǲ�
�+���hP��c����V�q`�(�$��)�,�_�y�yjh�:'�C������D�sHY���'R�h�=��݋��R�sՕ�oO��� �؉4E� KC���T��v���.0+ _����1�����>Q�3���C��wZZe�.>q(g��dq3mu�#�5��O���/U���Q�+w��5���ʵ��>�ǥR��(��hKN����ڱ���W�׺f?�t����ʪ������!�"�-���xU�$Ov�t%�8�; �-�q�}ˁ�\OE�:��G��e��A��r^z�Q���k'��Υ���b�cD�H��B}��_�Xnƣ��:UZ�k����	<��t���K������8���/3��g�O�/�磄0z�N�./�XB��f��	���3�8U$��;hk~��#�j[���8� -���+ɍԙ�]ڍG?G�N5�~���Rf��`Y�~���%���d��F:�wMI
lί���q�Z#[4<�L�}�7�m���7��NHI���q���Pn�/��4Q��DĽ��]X���f�!*G�F�$�r�k��S�ae�c�3�^�d�z���u��~[�?��ck`��QS�i��~�cP� �P�(�U5�֛�Rd��Vf�ӈ�Nr�����(7�g��U���.)����(r��B~�=Ζ5�� �ټ��CT�������x����{��'n�o�Qȍ�fN�=�T��y8�h"�c��O�m<J&-�I���PK�`��  �	  PK  ў,J               186.vec��ˍq���}86���cf�]�Cٲ�&�l�V6�d�M6�d�G�ץ��ק����>Y��<9�_��S��T�rʢJ����jT�%Ԥ���
Q׮��>hH#ӄ�4K�hn��]JKZњ6���m:hG:љ.t����DO�^����/��� 2��a(�(c8#�(F3���c<���b�Nf
S��tf0�Y��l��\�1�,d��,��R����d�Y�������l`#���Kmѭlc{1���]�����>�
q@r���opL�s�椞�4g8˹���z���B\��\�*׸nsCor����.��������<�)�x�^ڼ�׼�g�V��|�S*�g��S|�[��Ώ,�O��_��)�PK�Kd�f  �  PK  ў,J               187.p�y<�i���/e�Q�a�!#�2M+��!ն3$Sʲ** b)S��Z]�FR��%T65��b�f�1eˑc�����g�����>}���|����}T2�@s��� B  T/@�� (����H$����8,�������K6��%��ƆT3�İ61��b�Xdc��L[��,��! ��aq��L
���ס��Q�#�� B�J
��u���� 
�#�(4��P�	@@(���0�:��0<|��	A� �D�@���9��hy6ї�?��,^���k�Ԙa����S�6�\\�n�=�xm����۴9p��A�;wEFE�ݷ?&��Ĥ�BQ��S�ϜM�Ȕ�\ʽ�w���ߕ�߬���w_����6�<��i���]ޭ�Q����|5<�vtl|��ɩY.���?r��\
C�r��}��08�
�ȉ�� P��Y�]R��-����߄YLgɍ�g�ޓ}ء�D���\� 
������	8�����Tum�Q��b�h�CadX+4I(�k;�㓯=a'���&�N勃����&�����⡡|4p�7*��K��_ܿ��y����E��#T�::w�{�3���<2�%l��!��X[a�z<b�&͐�����𞸾��G������������w�SO\���S�+i銗JraĒ5�-�d����� �����g���E�/��fq�Z�6�~@��Ų��Dm:�>������^�)��<c�ΰ*�*^�7�6wՈK���~�ID��z�ɏ�h�@�C�7��N^��},Dg��ۭ��b�7+�f

�󮆴�[���%*g��.�Ð$̥U*`	�A�^o�Ǒ�)�S��>�pϻV�IOv�O�Q��2=[�Y�0��G�p��������RT5�4=]kDa0�{UO�s�/F�*�Y�d�Mϫe(�D��wu��8w)�q�-��Uؗ��%T�fBd0�p$�F�O�>�$Y�Vr��rF�E�c,�)}_�m��u�ȗ��>�D���z�<U@�W���}��3�De�3ߧ�ۋz��'Hjt8��;�ߩ�[�
�̦!�9�^g<��.K"b D�#9�B3�K{N
x���M'7
{R�4�~$$T�E�%7_7]j��Ӛ����>IM�!��"��{�6k����	1�@��;o�?�V{9S��Tmm.��!��n�3VBN�x{��:�M*��h@�;XbēK�{�g@eE]sǊ��\��!bd��odd7��豧�@�Ӧ�Q�z0f~[����b@���0^�p�Y��H�8\�ʆP\�`7�%"�|&���oכJ�u{y�e��]mft���)d/Z%�24r&]K���ܲ�FivCY�cFX��y�N�M�~��c�=q��J�!�|�/4w���u���)���S>�����u���ݗ~ڃ��1��ӻ�������x��%���;�-Tz��-e��c+���zԷ<��Hh����;X�����N��
���y�:yf]�4�/԰���Z�/w���*oR�l�v�3֥)m���^v-K�J?�j���X?W޵۟\�����5��OƟ�]��3���U��y���LbJ6��0�*��1r��^{B���v���W��ʬ�c\n�������4�OTm�PKi9� �  m	  PK  ў,J               187.vec�g�Lq������{ｷD����e����D'�Ub��D�C��w������~1gNDV�O�
T��7��L��,����S��Ԣ6u�K����v�iDc�Дf4�E�EK�V�ִ�-�hO:�ɮ�]wW�ѝ�����D_�~��` ���2��`$���2��L`"����2-�b��`&����2��Y.�B��%,e�Y�E��U�fkY�zob�n��c���-��m6�u;�����=�e�9�A��qX�p�c�������=�9�s��� .�e�x�W�׹�Mn���;�p�R�q�<�y�e<�	Oy�s��B_ڼ�׼�-�x�>�ɳ~N��%�����"�w~d)~�}�ܿS�PKX}��k  �  PK  ў,J               188.p�k4�y�����ո35;H��d��Qى�r���du*iّ��l1�d��,�l�&$�E5+Y)�t��KQ.vt��fcw���;�W�s�������m�}h�9�s@ ���>�h$�D�Q(�VQū�b��_hik��H�K�H��K)�˖��uu�6�M-,�������1�ͭ��sK@��U%�����]�� �.@�! Á����"�O�^ �#�(4F�(�` ���+���> �!�,����(C�~$�"��Pt���4L�
��Ǩ,ZL��dd�����zÆi�r������:7�M��}|9~�!;v�rw�E�?p0�P��	���8)�����f�����{)/���ZqI�������~��[{���aˣǭm�]�/�=�z��Fލ���0>195��G�-N���!8j��E���K��=���mH?��;�\,��![y�"�TQ���F��>��3���D�'�_\�**̓p ����x������%~������� U�k�����~�Y��V�Ɖ����h��y��.�a�^�<4�`w;PL7���8eG�W�e��v��F���(s#���h2��R{]��MXN}��>�`Ǽ���&�U��~��p�%�^t����+Q[��[N����y�z�N��f��T�-�@A�QȞ�I�㷏(h�*���^88�P�=��}Q?w��}�G���rcg,L@��Q���>�U|e[G~�`<x��.��T+�'�[�=5�S�j{)�Y|�n���0��٠�X`G���Z�X��w��T"����H��\&���F�^����:�e"q�]�e��O4,`����Mb�G���,�u :f{7&_��fT�M�$u�iߧq7viɫ<�ђ=}�̴��a�fI�<���B{/� ��;TRI�Q>f���ف,���pÙ��x|R�����VឞUr:[ m:[�[�K�M�)��_zTXN����y\q��&|=nD�4#�qN���V=A_��(����J�pgDO���RKJ�DU�zS��9Gm�T��t�&�-�'!�X��S��>��F�6�wS�S(�^��v��ȗY�I�W�e��׋�?��!�Ge��8�w�T��B���)m���7���J�\�%T��ViW�h �s��&��T�Ȱ��%���	?L��&�+ϗ�9�l�q�/�B1�{nKD��dwe�g'��4����e��L�n�ׄ���aח(�րg��;�7�����w�Č��"����%P�c��ؑ���:ꎆbB�	㈮�iZ��뿪:�+�>����Qf�j�P���_�y��^Kz�c![��Q'�gX0_h��[�}O1�3�Hl�+����ׯ�N��<74sO�PO+��ǞOur�����ha��e��S/g��D�A�7r՛�rZ�yE��j���o�Y�N7p%N�z7�l�\��I��'�����
��Bc�j��
��ƚ�C2IX�_
6r|y3�4�F��3Gz�������2?�Gp�)��ll"��N��Q[�$.�\�F�$�|��dy��k��X�8A,X��g;��$��\��9B��/�L���йR}��Q�������E���>����4�Z���;S*�RC�L�G�٦�
���}ӈ�������Sn��eͶ�PKD�ː�  n	  PK  ў,J               188.vec���q���>���ݵi�6�4ӌ�ܴM3�4?1�4��Q�������׃σ{�#�2�����%O9�S��)�JY>*��P�jT�5�E�T�:vu���O҈�4�i�E3������iC[��ޮ�]Gw':Ӆ�t�;=��D/���>����@1�!e��HF1�1�e��D&19����4�3���b6s�,��<泀�,b�y�.�Y��Y�JV��5�e]V��Z�6���la+���v����a/��ρB!�!s�s�c��q=�I�Sz�3���S>.�E.q�+\�׹asSoq�;�r�{���C}�c��g<�/m^�k����[}�{>�O)��T�/��P�o��;?�?}�ܿS�PK5�"�f  �  PK  ў,J               189.p�iT�g���C Y�!�%�B �B�VlX�b	��SA8ل�`@�f1D�%��	�eeqEİTD���L��t��ؙ�s��|�������9�zP�X�ś��Z  j�<$��Ð�Bj���h����>��������r���\G��H.v�68R�T���׮�MNT���B�u�ƺ���@��K}� A@--���6 ��'�T�?Ԃ@ap����[h���A��n��@10��f�!'a��R��J�DF����n�X9��������Z�ؒ���4W���^Lo�{�@�������G��y J����#	��i��3��y����HΕ��P^�s啚ں�2y}CKk[{Gg׍�;w��00��btl|�r���ٹ7o߽�_X����_��0.-(E,s�Z��(��7��A��-)ǐX����W��of5��mm#+��zv��K���~�7�# 5�A0 ��&IN��������.LF]��0�WX��+~�k9��a����^�^�IS�#�3������ڲ_0!��UX�\K�oA����X��8�X�Vt�&����}�G������{b]�����@#�[��.�$�Ӕ����5N��
v/|��ǺV��H�+����ښ���,\�Ej �@O������=+�3A�J�o����=>�#];&�_�����.��ht�A���.x���`Ib��H�/��ճ,a�]�~�u�G�܍�;�Z�ֲ�J5�<��4��(%ES�'�B���s�~�z��@�q��������~�����=6M�)�6�z/�����N8�׌a�ZK��XXIq͎��/����@�����J-=���mF��D�.���7q,�A��f<�$JЕUV�^��<'%�/D��eÙ�ʬs�$zIR�e�^������G!N~}�M�����U�9SO겋|ݵ{��c"��"�g?��Q���9�S���_��W�q`S�OE�E��B!��I�$��v)���oy�v}ÜXp�(�%�U�VO����4~�۱�����+�6�~28j���i�>O���o�d5p�E�W�1�P7H�h�>s��o)/ӫk��b���b`��>�Vc����;���[�X�J��=KeÛ���.ȝ˂]ߍ�X��F�+$/=�o��v;�����ǒ�������D���g����ǿn�.Z�6#w8���Tw\����O&JH�c_2�<NnkJ讴��*��7U��ҍo&�Is��.=�CHk���5�~���z]��w&XA��ׁ���~躖�#[HPU%̌>�ׄ�N�s|(��� ��1U�;��=Cg|]G3�D<M�/�`�';��fG�H��Y���������_��q[�~)q����x#�b��hMF+�y�rԑ�[Q�͢�]��yS��M!�H�I��P��|��V��l�������lng���� �����u⛤;�7�co91�a�f{7��~̚�����i���Ic����=y6f�WXN��FRӜͨ^��c���V�G�ї�s�G�&Ӣ���鰜�z���Ld�KS�\ʢf�@�y��D�a��Z���Yӕ���8�,�`��;�b�0))_�et6�����8ѱ��s���"�R�G�k���7dw�B����+r���n��`２�t@���/��<�x�t�������2W�!^��PKR	iu�  �	  PK  ў,J               189.vec�e�Ta��g�g����.0�
�؊��
�`�b+�b+�b+���q����zn��Dd%�yr����<�@E*�,*g���J5�S��Ԣ6uR!���sקiDc�Дf)��Z�[Ҋִ�-�hO��h��ݙ.t���AOz���ۮ��/��� 2��a(�N)#�(F3���c<��$&g���S��tf0�Y�f��\��|��E,f	K�,��rV��U�fkY�z6��Mlf[��vv�ة�������(��0G8�1�พ��)=��r��)�"����r��ܰ������r��<��#}�����%�l^�ޖd�N��|�sJ�%�k���R|�?����/����?)�PK�O��d  �  PK  ў,J               190.i��eTL��,��%P���@��E[ܡH��
ܵH�@)���Z��U��@��w֑?�ǽ��5��^��Y3��3�K�� rey%y   >��*@�������@���T$�DD�t��Ȩ��L��̬���,<aN>��� �]TB&��/ �w 11-		-�)�S���� �@)@>6��EĦ ������� �% 6.����!������������y�<�8��O��x���A,nT���|�LM7���/V~�P��4�t�l��98���ED�d_��+(*)����604�������w�x�������1<"�STtbRrJjZzF��¢�diY��ں��Ʀ斞޾����ᑙٹ��ť啭��;�{��G���/.���B_��`�[�G.�.,lп\@,�(pp�B�(��@�n�X`!�T2	5�~�_��ӄ�Y��~����d�w`��_d���\+ bl���aS ��_@%9*`��Rؘ�s�k �t�{��#�S������m#�%4<���iA��3H��3��f�m�҉�FhC�\�U�@c�%��	���9�8;~w�����D�r5��K6&j�Ma7Su2Z�ZR��!U�^w���!�J�'%q��q��mBB��V}��v_��QS>Y��&���E���;���f��v�]��q��b�$l�VA��*����f�ů��^�t[�L�X\���l�D;��c� �~l�d']h���ph����)���i���L4��p����l�NA\���-ς��5i���Ӵ��+?ik��A�l�)��uO�p~-��eԵ嵎����<A*���8<e�$��i6��*��v�F\�\����ƻvy�*�o!
ɪH��8�Y/TE�	;EEN}Y�kss\��E�/��BО�l�o��qym+l.o���w�g��������dZo��X�* ��s
J]��h�'���[�!J�?�0\���d@�S'Of��Y汇3)�%�|��F����R�/��gA�!�x��_��m��o9vn��������U[$o6,��"�SG~�o�����E�ϊ��%��L�1��W_�0M�l�g�<O>(��v}��S,u�L,3s�����m$%�k��q���d��)�3W�a����#R2��0:\l �Ѭ��I�]}�U��j2\h�D�K�΄���]ȸ��Le�H���0�WЛy5l��3bE�z����P�}�����qgs"��^��!̶Px+��nXۀL�N�d���D��1��RWnG���(m�z)~��E*ZX�[(I�d��Z���z�R������l��Q��O��.ެ"�嵎�"�==Ü�7�dWS4�ޝ�4ъ8[�����xU��/��`m��!:DG�-c�+�r3��\������.�ԓlQ4s�pr�'��oXi�Z@O�s��We|�O;�[�����zv�S�I|	�ӟ����?�ue�	z:/+;P͙eb�5��l�^Qd�^���#���u`�����]و�����8^*��z�"�Юzr1DXV��ū��>�Ã'�����s����|ρ�fD�C�İ�fk�D�����7-ܻ$�+Coax?�r�@���n�I��Q� ���:��V+�ĕ��+O8j)x�uر�~�2�qu��\����6����qj��qӝ6|z�eN���t<i�=#����>���A���y
�ĶI.�,�i���'�A�&.��7;zj\:��[��A��w�F�O��z�!5�ndA.���Rd��gy==�6��92�.���)�=�|��B
�V�3�Ӽ����*�����
���%���Vj�2�=�zY���%��\���*��!�5"-2��%h �U��F-=Y�4��.���8��
lrl���}��G	���޵Y� �����G(g�U��`�A�\��@j�Z�Ǟ��v�������3�"G7��<�*Y�J��<͐B�0�����%b�]�A0�ލ��1�m���H�tI���V��Sz`�����0�>]�|�bޢ%�=��>ozG�� � Qz���3̄����-6F:�߱�͏-�g�Ll�=�l=�-�xO�<:ؓ�旅�C�]�q��S�����s��el��*n[�w�*m�Bk2U�������צ��s,� U�������H�Z�����$�y�V�QF_؏P����	ٳ��/S�(�����6
^>ma^"Y��~�9f�wZ��l70���"?������l�RT���f��iMϻ�";6j�@{�Hja��z\�s��U{��x,[�P��l�G�.Pzm6؎�vnL�,�?��w����(�fpx2���.P�,�D�/̻��8�4*"�����^Pbpl�K ;�o`�%1@�%֟����}4����K� 57��0S�Hߎ	�g�qȿ�BZ�r%~++�p����[}�ݹ�L�>��OsҖ <i���pX��}oI��ն:�w��O��T�=E�N�)�F�@s��1͆W���]��*t$�G��!aFBN(�{@���B@m�4R��	���5hҡ�D��8$���S�F��]��V�~KZR:�`���c�?X�`J��P�SIII���N�(UyI2�
"���`�J"A�w㈞j�D�E��m��Ht`NE^U�iLݹ@0��ހį �������nl��1�w�w�����j���J�#��P<@�\/v?�u��>�N3���^���S:�T�AʐK���L��@l��dk�a�|�BP��e�U��k.u%�5a��%1L��6����gK��:˾�j/��9���2��^@�"bH5�.�7Kna��8��JM#��U.Or(i�$���JwY�I|ITb{�Vݮ�%���8x���B���h.�[�+�� ��=k���k���yj�����.1}W���'!Qv�oL�Dw��$��q����RNSIr��3v�����V��6*ND'�� T�Y�IῒS�nҲ���z����mT����Yk1Ʋ�>�����X�_�=�w*o��ܔ���f�O�>�Ϫ& ���X��^{��w3�(������9����$+rg%c��0��8�w�g��y�~�w����j~~�����"��/�ގ��\�x��_�Kv�m֮m���{,�����~.����m�]E�$u�{�K��%����T�� �j�3i�:ֹ֫{��OȾ	Q}��n��A�� TT��[Z�D���7��n$��8�@@E�T��ͣ�O�??���߅f-i�N+�:R�spp��8�WG�`����4S_�6��_��ŞyROB�:�/,IGfmD�L�hQ&53���@	��1����ݗr��<_���Nm���{�h߿���\���j�#}B79�5#�����4jkIz�N�I8�d=�~o�w�9G��(�60�1��/8NXaW"<�V77�E%s�@��,H��-��c
�	�g��r	�|9�
�����Q2�����bdǯ�w����b���D�Y�a ��lW�HƎ����W�jXZ}?r���^/c^<�����	F�zFM�������~3��.v2Qu�����x�N��\L2r �ʫ�p�Z�>�DK^On.66p���6@#���3\��4�y�%d�ш�:HYN���R�����-'φSlH*w�E7/0�L��=$O�l!�P�sa ��g��iHek�j����jۤ�����"�l���/�W{��}䢣M�f��/�lgH�m�P��%��s@$���s7n��M�s�*@�e6?�ZL���	.A�w�FK?<�����k==M�uV�<P7�*�^�@d��^��h/�:8��;�bS
�P)�?��A���~���*X��@�\�u(ۀ�@�����R�Mr���8�m�����Z�h�V�������w�_�X׸�����2�xM�?V��ےBGb9��\\��񁯃���k.(Y�Yǘ�ѺÌ1��Ɍ��U7}��+U�)�#�NqJU���"'&��I����+��ֵ����hDO�gh%� %��kHxLwf�ad��ؗPH�5"H<��%����p`��c��V8�*��7=��qJ�u�FҙqH���ˣ������\��	W�<�ˁ�S��|��Y�����9�e��"�]��:0���:�k'w��zr�7R��aLJ*�r\�~w�'�r�MJ�eR����pkv��wIJ|VGa�H�aC��N�� c��X$�d<O0�!�-Sq�M�.oxŢ�3�.�Q2_
t�ָ�ۊ��З5���^͕�t�kyB�C���Gb>�<$�Z�����Vrv.�zI?j!VK*,E�֋�D���(hw��-Dh�|Ku���A5��_� ?5L�b�.v�󬕌2k�lo�vPyQ���7����i��d��Ʀ$+6!�$����|>n]S��2�t^%�OudY�*r�M��g�g�ĭ�U6�h;䪁�A�f�jZ�%����B�M�}_�w��K��yeQ'��j�#AR���X�c%op�7�(� 	DM���h�^���7=�;�TVq���X��s�(�=���X�Q�/u	N��j)Օ�en�.�$슠�{�!1���F�w�n�3E��swB�N��۰UBz��|1x�:��K��B}'��8+��*��!�pѐ�ʛ(���Zus	����A����半7Z<YP�;.m�A���e.��>P�#���5��l\��p�_�wt�>��L�,��-g�,[���̎t(|�й��-�$ `:c�@I����ٸ7x�)��Y��Ӊ��%�)�UH���Ի�ŗã#�=iW�ĆCku����e�qz�ҩ���_bE�U�A�t��y�ےީ	���@�n/��WL^�^���׫^��KjFQRZ[�������o�mR9p�d�S(~�����A�c-:k=�	���ue��W|�.$u�;/3,�#�s/����F��-\bg��k�ݺ��Cw�)m�*b[\M���y-� ��Hߩ��Z�m�����U^'/��R��j�ҚC@�R�F��7A�<�i�T��܌.�f��Ѥ���H=^
�r�W}͵��z��v�;����
�Ƽ���i�g���r�#���&�p�5��P.~�%���b���Z?	�t�غ~-Q�t�n8��n��Z�/�j��_+���ݜ���h�p���ؖ�SL���U�B���⎔�Q�;���
qz��ޱڜ���@���g�O���Sy�Y�VsU}��iTD)�w[r�:�;%4}��x�z��Y�o�G]u�8�[H�O�\����xN�ι�U�}���8�d���JtF�[�� �f�\9��.J|H�^Ր��.kv3����s��(5K��D\K�PA��U�G���F��c�pW��S^��bo��ię��>@_����C�԰^_~��D�.%d�k5m38�*��W�=�U i\���1��~�XY���"�ŧ�W��9N�P{����T� ׵X��SM��[����@kp��R��~���y���\���0v�MuL`}�̷%�ўgѷXp��詒��@����<�j��ZRV+(�9u���0�.R�4��������x�f�8�-��[}C�,3�X�nJcpD���¨٦]f����!q~�����H�ȚM(��]��/� '��̮a�q0xr|�	S@�$f�p�T�AS �f�]��e5鰘��̝�N��*1S~b�9__�,�5���DV[�y^z8�q(�Y���6~��I��P�6O(H_T��J%[N��܊r^�.��~��!cp��ƻJ�`O}AWY���sa0R'(�9�m��%������y:OWb���[*F����W�S���ãǯ��y/ˠ�1�f/9�kp<)o�+�{��a?7�ql����n��S�DMժ���K���>����0��NY���y�p��� e���%��UH�6%�T�_����"uaumC	q"w��H�X�U��v����H��z�mW���{�Ʊ��1.��TO�J([�lVJɕ�z��+���"����n����r�U�p��Y�ZK���n�K^q�xW��41ڳ��Y������e�m�E��h7���dď7/��d]bC�Ă�-Lw�YȎ��+Z�k����y_�/y�6M�!��"����:�^l�~Nl��(]q���qk�����B?R�Z.v,C���,�x��G�F���ek���x��i�I����A�$ý�}fM�����+��������T�ֻ7�����ik���*X�5�婝�Ϛ��J���?٘/>_�翵_2U��vO������BC�9������_j��$��*� '�t�^~'9Qq�YV�; �c_kv
V�S ί����	4�+����E}eO��$#E��3Uܾ  �g�"l�{�k�f�����L�Y=�&ۄT���ة�S.�[Q�h\�&A�ToX�J<_6���f�74t�/�}������M6F��,4@H� #�n���XL�p)�xvk�@�d�sw"�̸�c�i�=�$����b���̋X%�m�9bk�F�'٤H�� ��B�w)}=V?��2n�('����8	�Fq�<�K;���NY-e�%㱓���nq9G���33�	��P�����W�5}4���b6�|��tؐ	xlF��Z���˚�k��6�t=�'"Z����V�b�H�Ia����>�+A��Q��c}߳נ]Qp��åIi��}�'��-���B[�,�I>�+���Zy�i�]`�g���r�&�f��:>���$��PI1U._���;LFVY6�4ٓbK�H�+�U�[���q-�Z#�d���͵��+�!�㔈|fqx(�֪MZQ(.P:��7L}Q+�2�[�KtuFv^�@X�i�p���wf1m�fk3�%��I~� M�T�$�T��Z�:�'Z�n�q{�B]z�.&ԠWr�X���(��� ,%�W�}})A�w�X�X<S�)}���{��LNƌ&\�!/�~����0��o���
ҹ��հ�VȌը��l|��]l���2?v2{���"U�v)�);��B��m6qn6�C��s��~n`�f��;�
ݳo�T�G��2O���H��˺z�o����|fo.����!Ё��L��l��O/�Ggր�c�2K����v�Vp��g��A.�7�=,���cvAk֗�$Z��ϫ��2��t��p׌R#�#!#�6-�끸"����O�nP|���}h������I���5�KL��&[�����rd���B��-Ch�H.K*�rb���O�5%k��v�^�Ōw�S����$FEx<|[˻��&UzB6��x�s�u?��1�L���#�L����r1S���Ϯ .]8w̟	��	�'��I9K�]o���R��ߊ��^��hЗ',E�Єco[6�f-�<i�K�[�X�/�N,�����$&q\h�}�!�`�	 �*~w����B���;�r�?ZR�{E�zcv�y_�f�u��X<1��R�8��H#X�,�! �t��ZW��p��y�<S�J�ɀ�'�g��,WO���2G	P�J���x��䠅+�8�}W�ǳ_�Fb���<�=1�X��pLvbc ��CG&a���,x�dI��0��|��	Կ�z�r�3��֬��yK�(Y�/��,��#HQಯ���"�&-]�K����r��-�x����cb�XV�Q/ٵ������T_P� �׏�p^�>悪��^0�c�ş�̮R�;���X��?'/��y��D����3���L�:��;]�	�!�p-���0� |���_e�:V6p��VF����f�C	`��ϧ	im�r�
����jZ���9Ts���9�K^4�8 �*���m�!�"Q��5xDֱ������������iɪē����N�g�U-��X���Lu�/�PKGO:  �  PK  ў,J               191.p��gT�i��7�PL!��� P@� dl�Hg�82��q@��!8қH�ʂ0�:��C�@$ �A3�3��ew?��9�O��{�߹Ͻ��`h�֖  Pp �`!H\�D�PB¢81QQiq	4NNF~��������@�T$�{�4w�P(yUCc��Zzݭ" 
�ŋ��u����,~� �P�@� �� y�=��G	�@apR%,"Hh� 
���p8&�F� '�!$�HRN7�Y"�h^�*iӿ�����ډ��QVQ%��S���504�8H�<deM���?������}��>������GDF}�p�b"#)9%��u凫�9���ʮ�WTVU�ݮo��Nc��_��w<�|�5084<2�����μ��{9����������w[\  ���ʅpA`0(��B"��08Q!nFGzI�t�p�̒�V���͒�gp���eR���G�/�������q@

����R�4#>�\����*ƒ�'�l�TI��W�C���ܑ�	
/r�\�EE_/����&ű�F�R��!Yt�H��;���mN���X��|@x�����q�F/�f��p�E��ԆR�7�eS�a�ޗ������X��{ց;a����bm��w�ա-����ɦ^S��"Y���2�Mj9�/"�1j�W�}JS��ɥ���>4f�̹��w5�3N���yE���F�j�fn�^�J�=�2?���ɻ#�܀���0y�d�b�]��4�t��~�>Р��]~ZW�X��-��ګQ\O���Sq�'r��
K/{�o�CF���l�Y1��~��57ˇ��IݾIQ����F��dU���0�\��Lݏ�'֛�,;�i��;򽍒�̟@}Ndn��S�rAK��,�����<!{����!6)��v�v�~�����n!a�X���5�U��q�-v۳�n��ˈs�~̻�=�ct۲�3�Ăx?��ѩ����\�w�ޞ���y�5w\�EO�ުh�`>ug[���y_
=�q�����$_~5���-;!VCwݓ;�u�,
 �z��ަz���x6��[�2/�q}�ۮ�'�vo�_N!��l�ʓ��u �v���G�������E����tSrH�k�A��J��a�K�#y�'��ZӘ�v�?��y��җ���5�k8��ʉ��t��� ������S�J��֔�U٭���.M!�0ԡ=a��O���3Wn�7���e�t��l���4S����nѸ�(���`�׈�)��O��;�[q:�5k��x<W�b����� ���yߛ�/mԂ�o������i$�+׺�$�r��:Y-�K����GG귂L�H�Wq\��+}���yP_9������A�!��d�o�j�/ݙ�̰���ۺ�T�	&��!�_ث�X#Ia*�H�������wR'����������5:���Qv}mߎy���hT%^Jv��=F	d��|�v=ej5r͕V6���z�]ߎ�(9W����u�q�C[��X=�Q�R�Z�k��t�I��/y�����C3��%n����6��rOx����NRCK���UɰU�p�|����9�-�	L��_�a�|�v�s��i��Xǭ2]_�O5р,v�/��R�b�2��W��]�S��NW�T�x#��p�R�Wg��6�Ϫ�����\N�4[�IS[���y� k�L4e��z:�A��|`�]���Z#fM�P��,n�7�
�p@ծ����q^ܯ�nQ�y��e�!������}���U��/��PKv�(�  �	  PK  ў,J               191.vec�U�a��5[?������l�[�l�l�Vl�Vl�Vl�Q���z�pͽ����J"����<*P�JTNYT�
Q�]��Ԡ&��M�<���w7�!�hL�Ҍ�6-�%�hM�Ҏ�t�͎v�ܝ�BW�ѝ��W*��v}�}�G0�AfC�pF0�Q�fc�x&0�ILf�oL�iLg3��l�07�b��gY�b���eYi,��d�Y�Zֱ�ld���V�����#v�n���}�� �<�a�p�cO%qBOr�洞�,�8υT��z��\�*׸�n������.������>�iV��9/x�+^ۼѷ�+d�^?�O|�KJ�5�ŷb���<~D���ʊ�����7�PKƗ��a  �  PK  ў,J               192.p��{<�������0c�ff&#�-f�0ª�6Q�uB�.ۺ_N�´!�Xjct\j��.2n�[d�QF3��(b�9�:��Q���������}=���|���
�O�}���  p}�1�@!H�
�D��(Y���è*��	jDM5uu���D��VW��o�74255%R��cS�M@4��è`�*�Z�Z�����
��!��p �� ��9e���!�eHZVn��Z���C22p�z5z��q2�ZF6<�I"�_.@i�*���KtL|�в�[UT�t)T�v=ӝf��.۽v�_8�sv9|����������'O����GDF�寉I�SR9�W�Ϻ���C.���ߊ�KJoݹ[U}������m���ή�G�C��#��&�S�E��so��/�_\�}y� ���\�u.��\ ,b���2B(ڰ��Ax�q<���\Pٌ�69$Q�	�U�1}�;��������/����k�@�zx�$]4nF���-�nɤ��q����^���3�*���*�����fu�c�A^F��� N���U/�S�qK��*`��͡v�~�ml_rݡ�k�o�_�Zc��������hh�;��W���"+������<���qo3�X��1��e��VѤ�߇���W��)����':�e��d'[���K$�������q�n������UzB���pH����1F>pW�J��3/�k��OyWt���~*�-��_5��x�Z��Z;?��i����U���AȲ*���{G)�6yM��Y�֚65�9�O��e-_t�ӵX6H��<4�D����#4<��WƬ�RsJh�S����_`(я_Ns9��4n�fޕ��(N'�e�2�$�s���f�0{Ҝ��o����яg?�����*pXX�����$�ml��M��������Z�?Ƞ�\��^y��^ރ�/��^*<~K��AV���L�Ƿ~�'�m�!>I��8�b�D�EV���'�]��֮�=�R )��Rߒ�X�wiם��eQ�Λb�\3Q���E�� <��Ξ���7^E=�Y��_+��@�[ԗ��b� ��>�]I�h'�3�h�yAGk�l=�Ig������rJ���:Ύ-nE������������ez����l;�A<Yr;2m��6����eWK��1�ea
g~
6���=�߄�m��\J�C@զZ��~y�\x��Bq�*��ş�ߞ����Q�;�U��T�?��D�cu������g�J0��i|X���"�£�d�΄>6l�k?��Z�����4.�҆#F%'CW�D��˺��~�{V����SW��������>o�y�^�J2��E�yY��@�M>E�&|�)�M�0�<�93�4iTy�$�Y���3��~��p�q�u��JA;&qg[�;Z��B<��
�RZ~s��Zç�W5�H�J��O��n,,�j��Ω���=,D,���+Y��yx��X�2}�y���t�3��97/�Z;�7b�*v�鄺�[����Wν{x�I��?��vKe}8�M��2�R�����L�.�wcS=��ԓ}:P��rh�L)^�>��c:��m�E�)wI
| �|H��sa�M4kp�S���>i/�~2u��b-{�LpS;sM�������(Qĭ�X���&,M~��jNd�h��  �fWf�%Ճ��ˮ���G���Y�#'ǒRg�%;��/!�;PK����  �	  PK  ў,J               192.vec��Ta������݅���*�b+�b+؂-؊�؊�؊�����������p���D�S��b�S��T�rʢ�]Uw5�S��Ԣ6u���gW�݀�4�1MhJ3�۴Ж��5mhK;��!��h��ݙ.t���AOz���v}�}�G0�AfC�pFP�HF1:+��8�3��Lb2S�☪Ә�f2���an1O糀�,b1KXʲ�,��
V��լa-�X�6���la�j�ng;��t7{��>�s��y��0G8�1��B�Г��9�g8�9�s!��E��e�p�k\�7mn�m�p�{��yd�X��Գ?���%�xm�F���|�#������T��S|/��G��ɯ�<~{�����PK��v+e  �  PK  ў,J               193.p��{8�����̘�jj�2�a�1a�1ÈQC�Rn����ccr���:G[�V;��`G=���ڮC��n\�*�RRT�9��\�9�s�����_k=��}�w�W> ��w�@%  �{��2\����H$���`�h���m�q��	;����D=c}��!	�'��P�t:A�amAc��ik�H$��PQѠ��uh�s����	u%,���f���~-��*A�0e8�B+��(���A���X�< �¶�PY��8�p�P-.C� �IT���3=ɋG���54��ܥO6����`n��ܻ�m��������=<��N��>s6������Ȩ�K	�I�)��2�
��sr���E).)���������jj��[Z�m�z}*�����īדSs�?�/|��yqi� �?��za^JP(
_��"�`�0��V��M����e�$H���w�'y=(5=��ι5��f��X��e�O�y��l�w����x>����:]l���sճ��h�D�2ϕ���>+o7����Y�~�.5Ap .��!Ə� S�om(�T�3iydqI��O~G ŲAO�.�*�RϏI�w�y�XO����o��<��I�bA�j���m��O���b͹ϚVc
���,y�q����T�%�[�������+�t�A�����74�6cŠ%�I�E0��?�]�2���T7hG0%�e>��Bxcqx��)�\'����4J�>�&P����,�&5��U�Pd���a�ѹ����Dmn��$�J��)E�ۓ��΂q��+�9�:��3c�e�<�}h�;�I�b���,̨ɡ;��m�L쨋����� DY8'�z�M߽ꈧW�J�Q�x�|J���#�n`���ɄQ�ˮb�;�Ѵu鲬�sҔfu��K%�ja#(/�cggn�EF����|�8~æ�[ӽ[JV�M�d�m�`n��i<�f����$�{�����I���,�}ү橧w�G;�UX%ʁD�s���}o�p�?M����[�g�R	�NS�Os�����<)n�\�����u���q��ӟ��6��]D�|�`���][��j��Ս����2nӲ8QBu(
0B�+zq��U��6�ϗ��a�Q�O�r����o復�pKūY{k�W_�p��rk���*�����笳�×�EA=U�+�]?�rnzƴy QQ{���*<ȱ��s
��_f��L W̼q8ͼ�߿,ڠ ���:֑�\�z��`ŷH%���A�kD�?���Лo;N�.�F0U���7X6)@�k7���pl!��w�ٹ��)	w�d��]�'s�!�M�~v��'���dܱb��_r/<еS��v��3R�A�z��27�H�Jl�H�v���b)v������Ck�3������+��x��Ѯm4lD�[�Ŵ0�b2%*�;-�h�拎/�뗷�r�z�mč�!���cE�F��ʓ+�`C���S!R���^���P�;�{]I���6�j���K!k�gL��I��vUL�o')�Bz�Ydhw%�|A�4���@b�b�%`=����C���6�ޭ8�����ڠX̐QU~tuB2K:#h�XJ_��<��G��(yJ\�w����E�D�ˑ�����*/��i��5V[mz^=-��WL��	��Ǉ_�&6�8IL�r���|T�J��`�vG��/��o�ŭf]��q�AegoH6�o��8�PK@b`�  �	  PK  ў,J               193.vec�e�a��g���݅���؊�؊�`�`+�b+�b+�b��~]2,����e���F�)PB9��R�
T�Rʢ�]wU�Q�Ԥ��cW׮��>hH#ӄ�4�i�-hI+Zӆ���}*F���Nt�]�Fwz�3��ˮ��}�G0�AfC�pF0�Q�β�c�x&0�ILfJVSuә�Lf1�9�͊1O糀�,b1KXʲ�,��
V��լa�/�N׳��lb3[��6����y1v�n���}�� �<�a�p�cO�8�'9esZ�p�s��B*��z��\�*׸�n������.������>�w��y�K^��捾����G>�/)��Tߊ)���)~��o��?�)�PK���d  �  PK  ў,J               194.p��{8�������f�i�qF�f8D�	q�!��M�v/���F3���P�F���ΐ�Q�S���;%��v�vۙ��\�9��y�s��|�Z�Y���k�K�/z`�-�,  ��D�s )&��#
���IJ��i�89������������J$R4��R���H�&�h�:�z��$ 
��@K�JJ�Ҕ�ʴ��DM 	 r��
 ��P,(jH�������@C Q����j �P
��`�ދ�~ ��K+SM�d�'*A8Z\jRլ�	ޡkFM�#8%��Y�Y]���K�����2,,YY;qrf=v���i/o�3gCΝ����}Bb�e6�����732���ݻ_\���G�����uO�[����w��������`p�����#�c��s�~]\Z^��(�w��\�u.�!6�@H�F W��I�2'�dThqH�Yj^������#�K|���yvm������+����k����̓b:0�#%?%�CɅ��N��+��h9�|��I�ñXv���a�]��U��˳�дsy��O�ƙ'�bz*���Kgvf=��b�&���������a{� 
~��7�L�	��F�b��:�� #����@Ќ�!�ZS��b�9`A�{��&�ue1���"ל�d��b���cn��sY��I�KE�Zzs���OLI�wnxF�JaK\f��-��z}���,�)��I?4�Д5�2���ū;��'����m�cġ�b��o��'�*����vuG���c���Đ��^��Z��J"Tu�Zw(�5�<��'xq(%[���;��Ymr�36��~;fא�az)���1���.0�EL����l��rG��Kѱ&8����l��w�+����C��ɦϫ&����rn�JѰS&��ȍ��]����L���m&N��D}����$ɟ�r#S������cQ�Q�^\�3��1	�s��cte����Y��Ԕ����9f)��0Ӯ�[��寶����Jd����D@�))ߙS�h7�7�:�/���k�jv=i���=#έC	���3�m" �0�Q�q������+���A�l��NU������:����Ǵ�
Xr���R�ځN��6�r��I������S*W�;U�="�F��*��=��f����*o�� �*���yY �Pb�Ϲ�ߝ��ݎM�YY��Y��]d�x}X��n�M��e��EA�=�3��Q�ó����t@_F�㵽�ԃ��\̙���l�����&���z~)7Y]����c�W��f�M�lI�˫���#�����[W�`�h�\۩��K,��-��0��
[�N���"�7��5T�o��q��XlEp$%?n��VV��y2��f�hրO#��Y�'6e�u7�J� ��ɪ_�}2Ԣ=��&�+M�T.Ou��/~�PE�;\0)Y;.�!͹��U9��Ѫ��+l��>�}�+�h2�.zG��Q��E��aW~�Y�R T����c�d�c2���x]2.��kO%Εd�r��)%�:5�	������+;��B��ͮ������k�ե�h�|��)�aH�R�*En���:瑭fc�[Z�Z܌��t�X�ʍ����2��J�>O���0�:�"���sf��̟��MWU��h����O���,F&~*d��!ǂ\��b�e��_�w�VjR�'y�,�?�/,�!m��o}�\�<K�Q���rֻ0��=vutm�ː��k#{�����&5I���e�ŝ][Wڬ&�PK�p`U	  �	  PK  ў,J               194.vec҇�Mq����cｲ�Φl�d�M6e+[�d�M6�d��u���K�W�_�~���:YId>������T�"�R��8W�թAMjQ�:vu��9קiDc�Дf6͵-iEk�Жv�Oe����s':Ӆ�t�;=�i�K{��S��~�g �`�0�ag#�b��a,��&2��Y1��T�1��d�����\��|��E,voKt��2]�
V��լa-�X�6���la+��Ύ�4v�.v����}��@��A=�a����K%q\Op�4�Sz�3���m.�E.q�+\�׹asSoq�;���y�C�G��'�<��3������W���oy�{>�O|N)�x'��M��s}�?��7�<~;�I�PK��:�g  �  PK  ў,J               195.i��eT�����Ѝ�H	�C�4H��݈�8�R�݃0Ā�4
H8���Jw� =�g�xs_�{�yy�:�|���{�3�Y(4��?�� �~�y@ �����@ BB"Rbbz*jrf03+� +�c��cA!QQQ0�����������"$$$!&�#%�fcb�L7@I�� �`�ؔX8�X�> |O<���6.>�����>������������Ž���p)�؄��l@�>4��)	 J��h�q���F=xHG�������WTL\BRJZ���3U5uC#cS3s;{G'gW�W����#߽�����KMK������-.A���W +>765��������G�OLNM����^^Y][�����9>9=C���������?���Eyυ�����v�(q�؄��@6>����4J)�BD�hm}=�]�<����߁E���/���� ���/% .�⸋H� ��^��_�~,����
[���b=z���̠� �j�C�Ò;�Hd��c��u}ҟ��vuU���R[98�Ug@��,/C��i����k�Yj9;]�� _���K����A��Y���DQ�y�%����j�C�����:����'k�yY��l��J�Ǵ�~#�`��'W��X82�������Z���C�����W<j;�>;a{�5}�wFU-����������|.t�?Y0Q�+Ѣ �j�s���Я��ƻ�F���`}�#�_�[A���W,�D�HI|��]�7ٸ�E��fw*��e���뺛*����UkwW�̫�B@�} P�C�(�ڛ���X�K0!0+.o~�S!��S���^�I��|x"%)�@���s;�5�P��L�_Y������趌`���AYj�i�ez��h�^��χ��t p��͈�|�'�CC�[)�0Pp3����<� ��������i�Z[|8w.�*?4����_������id����DR��YU�e@��c�9��m�U��j�����1�u�A[���K��<N����bt��L����d��[<��%2�(��}&I�$�o}�eu>MxY�NE�G��f�w��4�FA�q1�޻��	��M-֭=�\rj�w���O�8��\�M���m�-�;k��뒅��ֈh��� ��h�������+��d���9gQ�,�I��r����U�/U�A~�A�D��f����5�%S[AD�ZHXK�vDf"��l��ŭmv;~�S���3u���Aa�k��*�d}C.������ن��Q���>��1����]�$t���63�]�������v�Ɓ����1ɡ���j�I��'�,�XWS1�V��(�J���r�Q�z:�y����tz�_`�W�U���ʅ-9T�Hu�G��?x����+:�m���֕Yz����59�����|=����Y+Jk�h��cթ��T���3�O��_���"��R��d��({HWz�z=Z��c� �S&�q�y��2���~I^ih����jj�C�Զ�oԾ!E<�~���3[���`��zB��׻�G�Kg����f��1�H|�wv��NBN����K����4��%F�ȍ��b����M�1���uOYxDK�çR��V^^�SG�}��9�:H�#�~�$�҃K �/^�m��o�[#P�|�P�F�z���Q{j��~��q���d<��2��E�v>7O��5I[b�uf��;��/ɖtHY&=������}�A����3��3$�R~��W�A�ھa���t��!D��)��޼���_-�ݔa���u��N�5�m��3�@��R�W�v�ORX������e�#�� �������1Xf��<[ԛ�ީo�vh�zgI~A�bX�u̓/)\�R��qӠo�~H�s�GB��?�nLHw3�N�����ՠZ�6)3���PGKw�w�{�q�QD}���%g�F5�ִY$�ᱏ�0�m���Vʦ�B�/��ti8��S�����|�2Oi�PrH.(����V�.{�xg���"��h�������f��;od���{<�{�%el,}�p:�;G�ﱩ��ƪ!`�t�5vV-�*��0�mH޺=�S��8�9i������l��aw���(PB�hmz�E�v֏z���Um��J��M܎�7�O╛�rۗ�PDߛ�S�s��K����1Od��m~�alK�X㘣Ү�z����g��0w� ݄M�b��Eq�0��'�L��j����F�7�	úӶ{�;���ۮ�l�ШA-~g2�@$䥞��Ƕ���N�f7�ky�n�ǿ��n�N(K�7h�qH����x�EN��cE��ú�[���V�e�'�{�v��jU�l�F�n�UH��d8��Z�0DB5�!Q��]$�~6nR"4]7�c?��H`j$y���No8'�Mؑ��]I,|W/�\g�D oh`lF��dŔ�_֣'���sqXל��w��*�u-�Q	�^�(�[Rf*N*� '��
�����+��p�a&r_��*�۸�f��"[tw��4��x����zN��yÛ��us�Zo�x5����f'�
�Zi�lQtT`]N�=0ܼ�-<�}y�ANxQ� �zȰ��4|�����=����������-�,���FO �Ρ:�F.�m9��h����mֿe Q�q����<9]���:���c�>�%�θӻR��F[���P��"��E��&���.-�5���Ū��Գ'�ɶ_� �n�Kxm�d�c�En~�9��j<�8�2�]�.�d����ݱ���7�uI|����wMT��Y�KX)� �䣐�Vq�C���o~ӵ.�.s��bp+����/m)�i��t��d^�L�ꍤ{4G����j���+V 6k=X�5�KS��������6o�mNa�����R��R�g�O�9<z�M��R�ˤH��8�<�`�s���/L�����?Pxץ�1�3�̿�-\d�F�^�4����ta���^j����4*~=����Ͻ7��*��;��_�(Qh9kL)H�5b3�mF���� yV��*��b)���������Φ|q�7{\١\)�%9yQ3_�Ģ�?�y0�bD��Z�+��~�r�zD�a���`�z5���15��-�-4���nH�b
�K�%�s=�gԪu�^���yo&�&FH��ߡ�*>��m��E�R�ɩ߿��;�S`�)C)e;tV<ң�.�ʇƅiMؚs����!yC	}��n���i����ݦ�A��[�-��Cb�j���Wg�_���������_�_�F�X㰩΄c�7�'��F�G���u-����XP0y�ʈ�Q����א�WL}b�E�����bƋ��J�f�ru~7�UJ��Ezg��
O��P[�M����-U:�	R�P����m>ܷ�\�'�6}�VV�֋�<��=�Y���iq��Lՙ�DEՊR2��,�V6�����R6�ɽ���I*��
�ۖ�-�Sg���+nK/��{H5�|\�i oC`���ou�ʄ�u���sd�7��h�"m��5T��-��2�m�,u����G��5�A����A�f�B�Q́b�͍�I�,	�=���ka���"Asyq��(�:C�حv��՚�yV���e[�/���LY�����^�/�YqA��ɭu\%�O�Hg�YJ�
�H��݌&n(��.�=H�ڮ��`ݵ,Ϊ'������\M >��������Kp����f�e
��ir2�_�%Ӕ̠�H���-��&ǉ���Òh�r��,��2�L:�����Е��J���������u���e.���;μa�]��j�\S�,���ȔH�h?��yJu�ܓ�|�ʧ����2����f[��v����[72�N/ˌ�	��F�z�@���������Q�3�{=t:��A��?)+���rB��y3�9��c�555���>��S3���j��Hr���Vد۝|�R��T~��j�����E>�k,+�����|[ųR����
IE;��}�p�d�0|�UXvD���͌��
�l��iw:=�����d��곡��q�B_ף:���QЂ^�/L��o��Iy�F�G�|z'��x_c}֔�a��˝i4�q�߸1�+�tw��1��6s�f��o�t�8�7'�~���&�^#Y�y�]�U7��>/�/?�l(�ؿP����~{�.c&<���w�%���x�f(@�Ŵ��"i�F�����sc��y��Z6<�)߃"�n��|b��p��U�mp�Ig�݌W#��lu��A\ ��b��V8��'�5ξ�ΰF�ؙ��\:�w3�]�(���y�@�\�iz����Wˬ�t�peTe�&<I����s�F�ü�|�O#X��	|P1 E��U�d�7H1���|�~iv�U��9�O�BH��N+�}��ei鼲���U��zJ˲UH
p{�c�c]����!<����Ю�39Ek��8�U8��VEc�,��,������w���L2U��mGn��br,����%�F���X�Ϗ��c�~�`O55�lg9Ka��;U9�u�j�ɏ���{�c����>���P���5��A��(~*[��qޛ��^�t�Q��[�!I�3�Q�;oT=��~ �WD������~X	�S�(h�z�]$d��X)Fd�� ��f�PݡRw����Q��H+��'bUn����?�>P��y����p�eTI^�뜤����Q1Ќ<���m��:�U�Q�k���tR�F^dS(��۫��7��
S]5����#_߲_���ʢ�����]eS�g:��n9`����(���77�'�>} \�wZ��L�ޅjc��*|XX2F>��_�D�~�>M@�[rcu�b/T!�Bi�&>��>je6o۷�Fc'��JZ�Ot� ��z�`A�u6��Zݟ�j9�ϳ��"q���#æg�iPM�8�7m���W�3��@hȅ��BK�y�K�x�#"�$�p��R����Ez=�c�>�8?��h�c�������Ԕ��:���ݕ!�*Y���l������ێ�qO⦕6�A�`�13v-������{����}сR�N�aQrj���%�[X�Ç����f��:ڼ!�ˣށ�Qv�C��&TC�����)$����q���+)�j�?���L��YH�T&'��8(Pz��/�Ub�sZ�<�	�g�~z��4��B�k��(�ٿ���i>hQO����c��h��5�<����x��4��}�.��9����%B�I7ZM���I0�����_)%Ѳێ��4�o��}^��E��,�AUg:��q��f7�+]���*׻&��!�o8R�3lo;���fʯx�Իqs�;P��&�%�؂����j��NeU\[G-�ƛ�4�\�\��:����E�0*�e������}]ɞ�RX�s?�yr�^�֘ՓSVI\��]�,U�Y]s�y�<s\+ޖ6ґ1�}E���|��s���g!:3��@��B{��R-���ޏ��,m�z�9�������-�#�S�P����T������[�?�g������[�f(7�m	Z��]bJ*�l�e���.�ё�L�`եa��=�f��巘
�f�f#P�1'uV��j��Ed�D�����^G��j�?���/\����<�Z�]�;i�5)߽�a�%	R�%֔����ėH�2�9}"6����[(<�߉tvN��"�{$��c��뿄4���U4/�f��Z�/d���'��I��qi
2'��M7�^���х� �aA)�a��Uv)�e<1�u�̃.ф��}���iN\���᣾!3d�j.�6!d3[���.������%Կt�a�������
wMnf�����o�|��a�J�/���T��r��o��2�#h�T��K���MD��e���%��ޜS(�J�80�f%��x8eJ��yL�|1���<]œ�sD��.�����EF22�������������ՌC/�]��{���87;�S��iÖ�6U/8�ΰ�>:�佋j8�{�y5�/RL�CF�UxYB���}̟�.�t�*�Bz*v^���:��Q.&rX�d��Ɉ��#�XC}ƾz�O�:�k���2ў�Qq��\�H�/,���}2�䗛���� ��-X����Gf��I ��v�_��9�^�Lp���+�)UOFJ���#L��T ��
D)x<���z�SX�;�����)봢��փn�.�|k�[n�W}S���}���ϏtԌe�܊|�w��-�^���G����>�\��\7�4����M֭�n �N�*��@�����g�&�?�o�=g� ���&72�Y&'|���3���U\疄��G~I�oxg�6�;"!x�8X�w�rq)�}Y^:�B:w���T�\�6������8^��V����rO����~%��gͻ�/eD	}����~�.,J��ޚ�j�hX�z��%��FZ�~֛gዻ	aE����$�{5/3їN��v���A%�w{~5��Ҥ//n+���0������� �`�-�� ��b�ziJ�/:}8q�_�Eޠ�S�E!����cM�����$�y�'~����~������Z���AZ�n�� t�sb?�����/�i�ǲ)n�61�2Z��P�?�:�������9o��q��̊���lhO�}�4�x��3��,Q�-��x���6}h�T�t��&=�Bn�!�]h�T��s����H�=>tnW@�t�$3��H�R\��تUV��Y��~�'���Mt�S���e��-�_�OM��7Lm���?�"h�ߨ�R��i>6�<w\~���dԟ�''rH�7�߮Qg��}[q)�t=-E�oW.��,!
P��U&��ݤ��J{o�?rj�d���}�F�
�ߘI�WY�!O���=}Q'�@��Ö���T��D�5x�
M}{��}e��S(��WK����n[���Qe'ef�C`e3�8�ʸ9ş�3���u�U�]Y ��r�4��k�RQ�ҽ���q2���`ݴ=(����u�|��E���~�To�wm����W���?P(o��|c�ŨHҼJ�=E����c}I)��:��M���1*����b+Vr��$���5���S��ka��R>�g�B�GҐ6x�F��W���h��If�&�޼2�^7����^ v6|��{��ll�O��H�~���{�������{�_��a��I�c,~�:~�)��쮸��`���|a�U����+Μ�	��$Ȳ�t��S։&\��1n�{Z����D��N�>dal�+��5���ڱ ��	��g�-�����P}��q��e[Ī����� ���p̾��}I�"��輚ok,�=x�&EJ���^������/a�+j���&f����9���Ȱ�QO�u�:]�#%�N�r������?�#w��!�ew��;)3Hwx����7 c�G|��<
#�k��wp�ݛ�ل���Ⴗ�	��q�����
W�[.�LA��X�co�R���F#��p&dW���#Ꝥ��"�~��U���{�Iu�`�=a�	�y�
��iw?���o��Yɾ��fJ{Ua?���&xu^�qLV�z�7�Bϱ�F��}�Y��2J����=����äW�t�s��*rY ����x4z
� �1Y��I�U/���v�	 $����(*K�\�W�C=���)-I�AOH�}?E�?�
��I��13L��Զ�bE� �w�������<;� msI+�.�Z/���W9��س����0��PK���  �  PK  ў,J               196.p��{4�Y���$(�T1�LT�%BeJ�N��V��v[L�9�T�^��t���Rf�v��x3(B<�v�uZ-���j٘��v�ݳg��|���s��|��{%c�)@�����d  $]�d8�a0Y.++�@���hy99y5�Êhu-MuFg���k��`����	$IK�lkM�1� �!y9yUU�F����	����`�. ��Q �В�
�5��H��d���4�Z	���20
�HwoH�
��C��3.�ꆣ��9�p����#���8߈$R娪���1}��!���5��S�Q�>w��}�~��������K��"�����1���)7S��9�����ݹ��������/�Ï�U�5�u�m�NQWw��44<2:6>����̛ٹ��k��6����e{��A�ꅒz�@ `��H�����@u0e
C�b�a]b"�S����p]=�1�T��^���j��%�Wf��� I�Fv�j�����?��?"�'�/�J�6r;��/��Վ���?lcYĎi�g'�|������������v6*�>�eP�B4�
�/[좿S�?{�(4x�Y�=��'�~�#}�W\���4��`|3��m<��>�X0�L�`�^���Em��P>�������L�����
��(�-qpjX�K�������;�9X;��b�T�ʭ;Y/h^��'#3�@Y�>�m+M97"��*��� ��%˵qI9!���;�r��~��s�HcQܺ��^L�y"��"#�e�]�uvSs5a,��'�c�|P՘���k�n�Tb��Oч+��'3=���2��������p�Щ+vtD/m|N�,������y�����S�a*=��੐6�壬�^@uTq�tx5�ۻ���\~��~�7�T�OG��gP����Uc�:��}��S{�$�EW�co�\^��p��?���<��I�=Am��;�돤-Ѷ2�T(Ͱ���+��x?d���d4�d�V�yB��ѳy��:��(-]���7����0�*KQ��O���%d�+lUlT0Ĺ�f�êAg^��Xd8h�wm���wnx'�7�v�[���̥�`��f���LrP���~��C8��рE�+�mX��B�>�(l��O���#w}�isg���
'н���SA[ӶN���O��3�&��e�N����闺��[L�9Db�He��T���t(�} ��
(����ĵ�6����>�����qVo��'���qG�f��:���-_?0��Æw�k	E��!�����ƹ��cN%���&�	m��/�h��R�-[[hCkݕD���;�6�z.1�a]������x��}���%�(�,�&�sv��>#~��s���}�u��ЌlJ���D�.�(�\�|� �Ik�J��;͠P�h�>�ƔV�6U�+[v��7���yCb#��A�a����wl����O.{���;�-�oE���x��ܺf�;  �)�R�{��̃�b>��U����uuE>@5*L\l��B9��M:��2�5kG+�7Xqu���}�D�'Cvn�i�V5��bH�B�n����n�-�ۛ�_��TB�m<Zxw,��p�'�_͈�_}�=p����J��ȇ�^�";bg]�R��1���&i`ix,�n�c�h��c�I�j��Ү�s��)5N8��@6=t6�̰;���V/��&sä�&�*Dc���� `5��Luz���%tƔ�6�	OpZ���"<Ң	|��Ae�d�/PK���  �	  PK  ў,J               196.vec�g�La��g�1z�-z��ItщNt���(�Nt�Nt�D':��Qc�k�d�z���#�|d>9J���'�De��,��UsW�5�Em�P�z)���҈�4�)�hN��ڊִ�-�hO:���ɮ��]�FwzГ^���}�G0�AfC�pF0�Q�fL���:��L`"�����L���`&����2/�b�.`!�X����[^�c�{%�X�ֲ��l`#�(e3[����t;;�Y(�.����~��O%q@r���(�8�	Nr�X��z����<R>.�%.s��\�:7�isKos��ܣ��<��#}̓|O��y�K^�������x����G>�9�����X�����?�B�J������?PK{:i`h  �  PK  ў,J               197.p��{8���?3c����`d��6�w�:�r?
�Zr�)j��h�Ѥ�bȥ}�m�����)�uk%�05kB�0;��=�s�s����|�����~?������dc���� T  P� �0�	()*�aJp8�PRF�� UT�[54���۰����M����8==�N3k;;;,��Ł���֎�~�@ �*H̖-����?�} ����P@�(�Xy�0� ~P�)�*����(@!0*Ϟ��(
�ad㮨7NA�J8����Y�h�y���f��x������;�<��}|w��<t8(8$4,��g��O|�z*�B=}&=����y�׊��3o��dUVݮ����S���Ʀ��-;x�:�?�~���Ǘ?�319%N�H���/|X�.-�{� �#��J� �B��u/P�����(j���R4��t%�GA�g{pV+��W�6�{�]����ٟ;�_��C�^C ��H�l7�u�<�P��D�߯.Y(V7 g�~�-��}g���%\V������'?L�����*~6�h������I"+�5zx̳���9ydw�����uK纤��8^r�a��2�㜜N��I�xV_d��‿��C�OWc\Տ\<����P�r@��X�G
�\���{�7A�	����*��n��
8`�u}W���9�VGY+�qTz�9���y[�s䐉R[`�
,�M�,�{F��-�%�]&%D*u�?�/NK��1î��촌�w��D���p7���F�8��������+��UB>7L*[`kI)�iߺ���6�����+�k��3��`2���������7k���~�[���P���\̮kk�<�kT_��F������
ÏL (�}�/D�Q����"��F̴�Ye��;�y�_p�U7k��P��?�VĤZ��q�ď���U���ȸ����aVm�7�� x��A0�U\��c�L/���H�?�j3���ZW=�*5X�/Jj�5�F��Ya��G$�3��;L݆*��f˃�~>�ϖ��Ds�����2�������،����m��/'��]�=�f2��v��x��$��m�7���zȬ��C(��sqj��#_%�}W{�u2��m��38=A��}�*2�\fp�((�N�K����^��r�x�c��~��%�vj�e���f�@��k�&j�#_����4��.��)�Opъ�X��1��Ww��hvu��0�,K>���/�%'R87���Ѐu�x�6s�*h�o(|�b~�%���&���v��\l��=�� 7�&�7�3���9hw�YK�E}��>�$�75�{�����\ma{D#D�5{�U�[�Si�mu|�&����I�I��>�!�����h�x-qD�Ww��,4�^u=Z��nR������	]�DhWtE����:�|ki��|@��l �����X����{��:<���~s|!�a�n�;�������JmSz`�Qi�n1�XN��J��ux��i�n�������cJ���+������Tذ7���8�|Zb���'�ְuu+Gs�^����Ԣ�-?4ݤLB�y9�������d��1�=_Z�{�uh����Ó�Oi�]s.����"������Y�W2k.&�]ʕ�������+�H�(ۢ���S)���r�����Ч1�B�I�2��ѱ�÷�{�>�����̾�~�*>�B�FC�4n-��|3p��J�˰�<TQ��M�JF��2@�h���S����T%�X�eJjbY8>���;�(d1<6�j�!�PKFv�U  �	  PK  ў,J               197.vec��ˍq���}8��+{ﲕ�d�M6ٔ�l��&�l��&�?��<_�NW�ϩ�/�ODV>2�����H*R��)�*Y1���Q�Ԥ��C�T�zv��hH#ӄ�4��MmI+Zӆ���=���h��ݙ.t���AOzћ>����@1�!e�A	#�B��ьa,��&2�f�Na*Ә�f2��Yst.�����,�Jc�.c9+X�*V{kt-�X�6���la+�؞�Cw����a�w�O�s���0G8ʱT��z��ey��Ӝ�,�8osA/r��\�*׸���z����.����<��<�)�x�^���뵾���x�~�>��)ŗT_K����=R��g�ǯ��o����PK�-�e  �  PK  ў,J               198.p��y4����b	��Q�P%b,E����:��v,�ii��R�&բ֪*D��ܶ�h�%ʵ4�%-ZQ���)�f��.��a�{���_�{��~��y^�@��wsvu@`  I ~
8H8�!
��Bce���h5E9������:�C06����pD��F&�d2Y���֒dclF&m_B�Phi����*I�K��%n0H�=P�0������0Ч�Q 0
�#�()iɁy �@�P�Jv�%� S�5=W�Bࣰ���J��Ý6%/�[�Yp4%�������ǀ��3����V֎NTg�C�n�>G����	=v��g�1�q�	������y!�;���¢⒫��﫪kص7����k�������QG'��qw��߇�GFc��3�/^�	�_-��{/Z�����ƶ���Y��#�C�(b���>���tM�
=AQ�xR�Wy��g��V)8�/�L O�l�}2�mb����_b����$<� oY�0����e�Kc����B������ԋ��g˽�8����_?������$p�\#>�Jd1����׳ߩf��^k��l�
/z��:6ǈԩ�����Z1��k�ߖ� o�J �|���Ռ��C@L���Ll�8�<�V:S�_�E(���P'��/�Ae�Z�P�u��Z�W;ʙ�O*�@���c{�1'�);�[A�x����9#�eL���4އ
���������r�>��EB�:�Km���0C+V!�ʻJ_�N���6,/���YiW�O$CY�Ϻ����_� E�����i��2�wJ�G���P�C���Ԥ�-�����V��� x8�OU��zR��������:��RR(̓��C�3�E/M��6�o[߽w�}���'a.vs�I��w*�(z� _�|�t��c���.����Ƶ�-D֭��{��8~�1�6ZCBr�/1L����a�,�ނ�^�_j ��oOv�rZ`aǵI{+d���ǆ���Ԩ�S�=�~���q�% <X�����b=@; �4�/�4Z!{�K�����7#[��)z(���oA֛������n�L���k�^�{=7���|�Z�=^�k�"��`$�G%�Ђk�lE��B��S,�����s�l.�!X23=;eONr����;vPM���� |���[�XWܔn�9�6?ìm���II���Ɇ/�Ǫ�:�0�r���BR��h� �[��c/4B��}_�d跼����L"���I� �,�O~�e�j=��t`Lʢ� �z���s�d��D�Xv�a&D�D��@I: �[��v����e��b��&����D�����'ꢳ��3������ge����
�.�X����Hǐ'������9u�paI�nY8���!|ʞ	������C���r������Nޤ�C{�!c(��&dE4��z�-"��)�O��"���2l���'k^���E}Q�A4B�%%�6��S|��R��������f:Z���\�Û#���UH��C����2��DVm�Iv Rɧ�|)�p��.2b���W�I���V���Kב�29���*���q���	B+�����x��AV��i����,2�{���[���9bqJ���&�6�ͬ��?��Nж��`�F-���ҏ
!s9�C�B��	m�M��+���>����m�8]�4��t`�ŗѓ�+Y��}7��d x�u��UrӪ�)[�c	a?��:�Ƹ3aF>�5���Yr��)�`����t���t)n$L-�k��l�y���ek����v��m��c� PK��	�  �	  PK  ў,J               198.vecч�Na���yx�W��e+��&�l�)[�d�M6�d�M6��K�������<ωȊ��
��<��T�"�����bWչթAMjQ�:�M��gW߹iDc�Дf4�i�-iEk�Жv��C��:9w�]�FwzГ^��}�G0�AfC�pFP��,�Q:�1�e��D&e���S��4�3���b���ѹ�c>X�"��b]���R]�rV��U��Y�kY��<���Mlf[���<���]�f{}�}��6��9�Q��b��,�㔞�g9�y�z�K\�
W��]����z����.����<��<��x��x�^�*�x�o��x��x�>��6_Ri|--�o~��H񃟑ǯ��o�?)�PK�z8�h  �  PK  ў,J               199.pՓgX�����L���CV��(e�԰®�aB�BQvd4&)
Q�� U�"P�,��	�m)3l�@/�����������yu�s��s��H$��ݜ\�  �t �׀ �B�QH4���`刻�de�T���ꪚ�jj{t({��騩A����LMM5)�-�mLL��61�����]��ZjZ��$M N���6 Áp(i4�}"���g�08�B�`���ջ��p$���&K���2�CAh�h�qZn���}e�±�E]��s����������55;`nai��Hwrvqu�<����{��
	=�q���ظ��Ĥ���ٗ8\ޗyW�]/�Q�/)-�����W�𠺦�N𰥵����:zz�^��FF��'&ES�3�K�+��[]{��p�_�_�pR/G���@X���e���1�A�m�4�}nqe3F��آB�n���鈞xK�w�?'��?��[�?^C��>ЀŇ?Id��?��X�q�ŝ��;�]�^�:��1�vE|WՐ�j��J^.w宆�j/��O3�7���~������`��	�
�Jg�u}�J��~����݃k*c�����<ޭ��(w��ݶ!v㹪���	l��)m�O�r����G��(��'�m\��p-�V�>�q~���O�[���,��դE�A+hl��`:�'�e�Ř+��y��S��G���l�;D/�y�=�_�#��q����҈z�< �ٰiw)�^��J�a��E-?��3d�0-?�z����zB7]��Ƞ����$�Q������.�i
���/ώ&�v[���l��3<��q�V�#�m&ĿD'�5��_�<=��ʦV��ިN7��=���	=��\W_F:�P`�Mv�q�2�'2<��<�8_���\|��j�;�^��o�&5��n�u*{hђ����,7�Q���ow� ���2�D`��ѴX��	�ycH�ڻ��RP*�@�7���GI"��0yg�����F���LoQk�Y��#{�7�H ������4D]0�I�&�Nan�1�yR-�bZؘ�����sa�r��H��M:���<���aB�o�^$�W�Z������F�����E�&tG+n/�)e�y{=�d��9��6��ؖ�]���l�d+�����ֈG:�{�7HS���<�;Ý.�n��f�iUmW�����I�����|������M��,�oP35gIj+|�S�+�\�)��t�����Ii�7i=��g�c�5Y}	�o�L8c���
Z�oI	H��d���R�)�I�������݉���|��zS��ǵ2�)��l3��r:k�dl�W���Tv_�|�����dN�;��4�;]����H����	���h����.*�<�-��1��|�cFoʔt������� t�����:Zt���\B^��M�+�Y�
�v]I�A�o�-~���!�ƻ%��R�iN0�j�^"u�we7Lxe/�W�2u�{�s�4���\�S��P.�1k>���}����ƴ��h@aC�H��yf�$nQͿ���=řm'��o]��S㬲3K���uZ���SҨ�^=�3��9�v{N�b�n��-����L�R ���lYQ��O�Z��D��N�"�0r��A��p5r�>���	6�eQ�'��P�GVc^��D:y̤�Y�b-"�z�W�Mckس����tu��\{r��\�5���]�2.�G(Nǒy�}�[6 M	��n͝���7L�v�J��PK�5��  �	  PK  ў,J               199.vec�g�Lq����Z���X��]���-��D��D':щNt����>��L���L�g�DdE��PH�S�jT�Fʢ�]-wm�P�zԧ)N�Ȯ��	MiFsZPBKZٵ�+u��-�hO:҉��O��uqw���AOzћ>����@1�!e��HF1��,�1:�q�g��d��L�iLg�d���E��y�gY�box�.��L�����b5kX�:ֳ!��F��f���mlgG.;u���^���������(�8��℞�T��i=�Y�q�6����U�q�ܴ�����]�q�<��c}�S�����=�}�;�S�>zw��sJ�%�7��M�"�w~D.~z�_��)�PK�<,�e  �  PK  ў,J               200.i��eX����Ii�Zr�XRB�T:����t�X�cQ�DAZI�RziIa�e���?7����9/�<�ϙ3�3s3w��7��� �p������������QP�SR3�PSQQ�32�1ss �rspq��K����qq	��IJ��� T� e	i�!������f��a�����. 9�����@�@@�@p� ��IB���F@HDLBJFNAIu��D $ ""$&"!!&����3�0ޓR'e�:���1�"S��4�Y�&����`Q��w��9�
	����Ƀ5��ut���-,����:�<{�����?�e`PpHh���ظ��	i�3����KJ��+*����[Z�ڿ������595=3;7�����������=>9=;�wq����� @D�?����p�EHLLDL�. �80�ܓ"eT��9�1�"ə5R�)��͎X�`���2�������d�w`Q�_d��s- ��n�G� � 0��n��R��f:�s������]��S�y��������������00U;gjl�"��a�G��������p����]�.��)}+�#t�.2��avޕʟ�G[x��rx���S��,����@fP��&%�0��p$�q�?1Zۍ��rh���{讏p��	9C���F@GJ���O�k��İ/82����ŵ��h��?��	f߄�K-�o�cے�7��!(���,�e���!wsg��A�o�:��}���"�M9V)�MI�e-`�����Љ}�R7d���vC��m��w����Q[$��k�Z��2�}&�Ϫ�ߔ�{�����蹔��1��e������=cG�S*� �$��b<o�>��!�Θ�Ш-m���O{BL�e=�8��~9��=d�љ�X�ea�^��p��(��]|���+��z�vI/�_�#�K>� 96����a�{���3����B���U{(+k�[:�ǝX ��e�V΅�:}���A�[�M� F � im��UR��
��z��:4�bz'�6|W5/����~��� ���H��a����:ȏ�����r/2��*i����J�
�$�����Ъ�,9U����=Q�t�33Qu}���X9{7_g>nuVox.�\k2/��nrFZzLH���GN�٣|�aH���7l��#�%;֧U������f��b�~|����oqz��\=Ժ�����R�t��a��dm�n����o�?Do���|��n���(f!]v{�VW-9b\,O���!��5[M�A
��{XM�h�R%-�Oj}�զ,JS���!"��36�c!�zD}�)����+���G�L�Z�}�uUe�OM�ք֣�p�1YWD]�c��_j�Lj��0[������è��L��5/?J6~���'�6e9�}?_�)�U':/.|P�r\�TQ���tg]t�u�$O��N��0�A��?�Ɉ_�ﵾ��;/��E�\gFk(5z�St�vEY�xRh���"DyYN�ĥ���Z�� [���<�N���R��Z�BU�O����+L�Y�=��J+祯�j����}SGy;�`���Ǟ���%-��u��CCC�4H�~u�g����{N`�Jpɀ�f���}�I�7l����5��q��}�*DM��Z� ���9��!���,�Fn 35�
Y2���l$��eg���ۅ�� N�Һ���ߔ��(��6	��d�O��jN��?���hyz��G��K�kv���]�y�~���9���s���@	��*�YAu�y���8����A�K:�I�BQ�e2���H�)MW�`�:�9��s����k��EoT�h�C��ܦMm�U~"�[�/O�=��X��	�V�l�?+���й�I�Ͷ��:Na�Qu����i����3ei�>C��DW�;X+����B�j9Y~QُC��O:�ff��;ə�!����/�6`rJ ��������8�:���iV�
_���<B^l���Y� �R��g1����*s�� \��������q�o�Z}o�}(b�6�i_�%Y�0�)�s���Z]C�}�������-�`��Z��z�K��1==�14�3���F��<�W�(6��s�D���f� �-�.����KxdY��D��n���v��<�D��������pD��P�q����[�z<�ɜ xܧm�P~��RL-R��+�VŴ��f��Cͣx�E��׳�+�y
���0�ك_m��f�l�.k�X�g�)v�̚���'Ϭ0�&��j�n�su�l1��EƱW���H�IHm/�p]� ��F��b%�N�p�%k�}�%l8b$��g��C��"Bȳ`@E�ƟI�<6�$CFh3�,��J�凉��������g�y�'>����$I�*��\RvV��<��wܓ�UZ���P��3�'@*"�Io`�1�.N�|K\^�WTԭ	�"����z��A �$���p^m����V�Lt'����z�!L�\�M� WٲI�[ޫzi��\��1�ֵ�q�F���L�`v����'b�g5Q�Z;�o&9hր�T6�X>���+B�k�/��T,p�f��R�b�{����괏�CZ�[wl�F�LR�y�ԟ&�R2�~U�߽~�H����b?fNP�o7�%'[Y�uDg���3>{@Z���o{yP�t�ok6��(���~4G�"�J�k*A�jyF�x��T�"�p:�����ю*��<���&笪�c���P�sP��82���i/}7�t4H&x*�5��jX��Wh����7=a� ��蹽�b�u-W�L�����=��C�r~?��ת� �$]�[��a��	IU��D�%��58J��e��$ g���I�i�cg"���k�q�[^�n�S��kҜ��3銂#ׂ:��G�X�����h�(��4m�)����k�x�7��引4]tsQXBR6rJ���'��^O-)��L��9h�K\�\�������/��C�A�۪�@n�D�@��e�����F�ˑw=�0�$�߲�v����o�j���A��^��Jc,_qUޝ��Ԧ94
/i��K���6��zT>�M�6�Mq�yZ��b52K�m�"�yܲڹ^�b���5�ln���M���H��J��Y=�7�չ����Nax�7�l�bX|l��R����˄��v�� 7b��������c\������?rW�L�g���Ε�ۥ~�4�"|Ɨj%���v�*:b�:�.-�
�_!��6�02M� �׳�U����g޼�3X��#�@�R 7�����~�栢Y1]��,Ӛ��4W�8�U�t ��U�O�[�� �N�`Y��	]	�dDUq
��Y��������7t�}k0[�TCd^	��2�����7�� �7j������@:'�e＋�]Ҥ�Xg`�H� <��� �;�U:�%��,PE��,XQ�*ںģ�0���֖'ŏ��,���/�?}����.'�Җ�:~� �X#���ZT�$�C�:?nh!���ɚ8�!����:�;���&�'Bs���k�ք���4����,�����,��0���{s%��&�C��.�Ne�t���osi5�?a#%�W~?��ʮz����~��n��Rm�{�s�=s�I+P���l��w�/�h�!3Ug�Vݟ��|Z5��x��;Q�-M�3~�*r�V(��&����[`����S���:��mjG&�D�.��J�kA�����d�G���}���.����1��^`U�wd�sx\�D����Zp��D���_|���	�����̊��{���$��ml�w�%ȧ�,��&P���!z��C9����}(����#H<d��|�S)P��DP����}��Z&���G����:�����9Ȣ+d�o�P�W����RtN� �����2{� "�v�G�W��9�����m|�?l}� ��<`�*�����s�+"k��|�8�^��w��ے��r
p�g>�R��~���{�/¶9�O_+�Z���Ǚ�)�:�#z�$�U�F�*U�e�� ��?�r�������z��2�W���U?7���o�����?�#wh�`~l��N�b��A�<�;-m��N���+��OǊ���~n{���S�q����sf�y�F��U��ܰ��-�ز��`�SFY��U�<�P����L�ة�nѽ��μ��:Z.P����r���0)7�Xn�㣍�y���瓚S����:��:NK.����>
+> �*i�Hb�\ֹV�&�V����{��8x:S�����o�m�Ѽw�H�1wt-d&�i�\ja�@n�9��_e��*^��v5{���ui�v�}ĸZ4y&"���'oߣ���Jk�U��p��\�}�t����P�~�k�'�|`Y�E=n��DrǯO~%m�?�M	rMT�W���oS�� Db�����I��Iԣ��o^jݺ)���Y�{K��r	��婻�l�"3[t��M.Z����swuwJ ���z�ŋ;�#̞z�B`��U�;G�}E�㯌���:�3�Xm�G����WN�:�Ň�2��/�B����V�Vm
}����3��m�O\����'�mDL�+�k��^.%DL�l��*Vfz��7?}9�����,�%�uV�Ij|Y�1u8�Bw9����Y��SM��������?dι��,�=�~~_��.���C5�6٥�ѿ�� `J_����
4�1�8������\桏m�$2�%7�l�O��w���ߩi�P��ܶ�N��f�g������,2;W�q����b�<���%�Y�vn��2JR W�<�Uq�'߂�����Iv�51�yg�j��,+r���t�h+�v��
���NS�d���t����	`e#�(�(@���a�
47D������'{TvᗦHg>na�b3����
vl�/����X�:�c�9�,��`�rm�e�L�	601��p[':.��P� #��f�4�����u�����:�4���a����k+5ʌ�/7�p�Ćc5�m�ն�	Ѷ�-b����kՆ��Y�M'�����>��X��ChAHb����O"t���u��}�9�s�c�Z잼c_��n�;�?�8����[�ss��+�wn c��O�&r0_>��BV���?iLh�����t�ڕ*E�iuV�=F%��!ґ}�̕����:�v-B�69��/���Mwk��a����Ah�1w���~i�jO�+����̵u<@��i~�z[o�O�h$����%J�bXլu��r�"���t���L��)�'�E����଀b�jAK��Y���U��15���R(��� �)E$�֐�	����b���\^~^H��KJ'����I���%��	�w�Ø�r�5(�����)���9�� �`�@M� �1]~�`IhցpL�;3^FM�R��~�{�id轼�O�HM��ػMD�ͱ�Tw�6ǁ��F|#���>��A��Ԧ�L��ŝ���Ǆ��s}��e��)��yM���ɗ��B6zʴ?��99N��r|�;�)��{c�����[��@�m>-ʒ_5Ͽ$_?�3��xZ�R�����d�\�����1�E_����.�F��i]���=�S�I��̦��/��&�~�:��.&p�)ɶ�s��a�[��Tula�hR'�V�����N����ί�%��/��CYK�x�~����8��3��c�Զ��C�~_��]oչ���#�7u�I�H��Bs��U�>�����I�I�S�ߜv�Nrތ��f�V�N5�v���/�7���],�se�a�#��Q�/Qocca������_^Y3"�����FO���e�5U&�86�
��ϭ�D^	ֱu��_&�����$?ֲ9OM+�7o��'Oq�X=�2p��t��X~;�:-#�0�m��/ �n�<f��PmfjឪI7]��ʐ�������,a�	sR&anP�@�nr�ul�h�3,��6:����C$7�P���Br��V1��n��?��G�޹LI�4�<�"�m7���|�tm8����k�~���ʥ{�o��R�ߏ�����E\,���4{��+%m>|�*�#;/ܧ.Tz�9`��M͑���r��-���O1�O�>G�c���� J��B��,�Ϯ��--��a�'�����rnf��ʸ�mK��v�����!Y|_�R�8�϶��<��g���4-�ސRs�Ǔ�ܝ혆���۷E` )�/T@Qn���f�?����1�����;�� �ԁ�N/O<�vpի���F�5������|;�cgUbq�*�s�������"��zS����SV
���%֓���
��rBw/p�4�y��A`�؎6�1E.��/���(�E��Lm��V��FAN`����kQ1�	_����n�?���s�����<|Ӧ-g%����L��&�O�(StKc��KB?xNx���U����!k�al�ؾ��F�}(�!�w�+�j%�2a�v�/j8���Yc� ղ��됍��O�{׊aQKi0eL�/Aw�x��u9�ct�Q9�τ��uZ�=}�q}5p ��KA�����M�epŗn/���_�9���ĉ����|!� _g� '��{�a#F�~5�������E�S�S�g��b��][�6Ku"g�H��|�q�3zq'��^�v�����P�ZLn����CKQ�5�px˺���w�9aXhZ�(����GS�ݣ�S.R&��$_�zE47�?.�v{%?��Ե����)���֎\�><���vM�ڧ��2�i���'��)4^۠2(�����ws�"��X?�n�;԰�C�6ϰ������i��6"1p�tB���]�Fxiyh�3uV���L`��R�D�ͳWd�����@��(A8��#|+y�!�иy�'���h�ye63u=c�.��;���+��[��`Q&Z���ϼ`�*����� ��n雭S7����e�� J�rW��"s��d�Z�Y�5�[�J��r��zR�/>��%D4��l��G�-H(��Ӿ.|#�b�Y ���IZ��IQ��D�� =9tr�� ���}��O��QCV�Dឺs~-�kV�x�c';�������7��6�Nk[l�ǎJ"V2��MM;�$@U&�C��i�ʱS�T�J��5a:���SL	�S��O�v�ʅ���}Z3�����R�*h�Iq���0��+� ��?f�r��A�&��Kx[h�w
e�Z~�m��r���p��3�B�^��$��淈滏3��� ~XMܹ邗� ��UL"�'�������j�Y%�j����Jg���ջ�AY\��� f�u�o�����x�?��gX��1�\?9��]
Bh���1l�NiO��Z 5�5o �K�q�w̓:1�z���?�Ym��:�ځQX�nMZ
�2@�Y\b�����Λc&t=yW�0N�d6KN�࠰3e��sr|�&>�+���h�U[�`�x�s��}/�e��>`����0�\������d�%1�wHAd��m|V5$&�k���+�ۺ�,���`Hz��jiO��|���oo��Vb��������U�����z8��f�9��qU���~mXj���u� ;��A5��L����c�b;�̫���O�۴g ���o I�M���b�ޖ
(�����.�7��RXY����m����,+�P4J�;J�Ջj�g�@�����D0��������ɍ��;z 9RR}��u�Ў�R����cS8J�s{���)z+��x�����L����Rϔǉ_
ox�퀔����h������f(v��f�� PK�W�}�  u  PK  ў,J               201.pՓiX�W��!�$$���I�eB#X��XF���@YdU�HX�0�CK�q����M, ���%P�������P-|f�2��|�s��ӹϽ���n�o���� � �$؞���TF�B�p�,#�D �*��P�*�SUW?@�'��%��SL��h4�~�(�L߈F�9�Ñ����2UC]��_�v'���,�r0H�B��h�v@���},���C�e�0�,B��� H��`)XZ�t�I� -��ah)��q���2�*`D��.���$���,��~%eU-m2��!�����c�6�v��N��q;���s�~��������r56.>%5-�zF&;�������K����s坻\^U�w����ֶG�=�}��G�2�Ø`|����3�s�oD?�]Y]�o�����`�?��r�%\R��I]�ـ�Hk�(Z2�"�iR�0�U^E}�htz{1��~�����d��"�'ؿ�~�`�dx`4`,�Q8������pڵU��`�$��4�WHES�t�����9%��Sl��S-��}5�4��Q8��k ����2Ks*ie06pJO6Ч,(�e�
F�0�b��R��������7��z=��-����N+�(��,�
�>�r�`�
�w7O]� N���������9�,�ԨM���%D�c�@��̸V�Z�����ՙC���_�xȘK�NjEϝ(�F��>�%�+������_�xg�M�,1���W�;4���X�Y~������u���W�M)�M�OzU���gfk�[��:sw��"TSp�[�/�rÜ��{[Y�Z!ʫj#����q�Ÿ!w���o���и�_C^��g����F��3?܈�k���n>�=�����]h"As��V�q��z�x�M����� ��<�PhIg��3LP�ĵ��� �X���=c�<�Χ�!%�b�M�4���)~��������ggu�ؙ�v�K>�%��z��O^�vn�ݜ��԰�v��fQ�̆�[b�S�ؑ�Fֽ��1R��fP�O���|��wT`?��6j��vǔ�g6�D��p2�I��۬�.�ؓ��g7y��_�7���Z�>"��f�u�B�-�
�����;�MO����j��JW�p��aKe�2X��X�7ڋ����_��?�hO:6&��.�hKH�<;�����l�^��MN�4�u�]T��eI��uR�������(���R8M
�k_�p^unVʥo�J&�g ��~'�JfݧG�Sz�ik��N�I�cBeK��"��X�xxBa��U���p�zP|�$��6���p2���ܺ�E��>�^k7�0"FQ���-�G�-	%f��\l�#�К�8����N�n:�u�类�I��Ue�wnҭ�+!���D��|�s���c�hR�3ܜ�鎭&�Vx���#�Pi
��{�e�#?0-��H���@��w��׻�V�o��6�%���RX��3ec^ESt���u�KG('�T�6�]6X2��q٤�]�L ]�l�!���J���9l
������״�>��b0ˬ[����i7����j=U)
Om�iQ�h�A[��"Z�����({|"f��7�J~��\����sb��6��+�="�#�9"uh �0��"��{�N݋&�;���:�e6n�G(:�����֚��T�����#��P�!�}Oo���:~{��q}����D�`V)��;��?��S�,~��X�]BM\��,6�E�t�-���*x�s������u�~�m@P�׺�[�ax���v��k�ᡖ��]�Z�|�v��5�L�L��bU��
���f&��Ϟvc.�{��ۖ�1lvK���� PK�0�R  
  PK  ў,J               201.vecч��q����ww�=�>��le+[g�:dS���M6�d�M6ᬲ�Q���C�=��z��W߈�(2O�
��KjRL��Em�:�ԣ>hH#S�r�Į���iAKZQJk�x_[�2w;�Ӂ�t�3]蚪�ܮ��;=�I/zӇ���?� 3��c8#�(F3��TdY���L`"����2�f��`&��d6s��<�����,b1KX�2�����b5kX�:ֳ��lb3[��m���`g>�t7{��>��� �l��r��HEqROq�3����E�Kz�+\�׹�Mn���;���y�C���>�y�Oy�s^�W��MJ�V���|uT�?�O|��׿)��R|�?������?)�PK�T�_`  �  PK  ў,J               202.p��y8�����1d�LɾF��uec���4�QƒH��M�&�j�C�A��xH�t*
I'�ʞ�(DCs��<w��^ν�}������|�����~���+~#dh�T{  �����- �#�0	�DJ��8)��$z;VvNI^EYI^QQ�`�������H4��34211QѶ�cN�m`lBZ��D"ђh9))9����?�} #�@@� �`@�V@e�O�� � 0
�#$�(ɵ�;2 ���
]�F��(�U3���ҏ!�O�H��6U�N�_ƞ�qH��mr��5���:;Lv���[�`kG��8PiΌC�]�0Y/o��~'BB�¹>>�BbR2/��~��k�?	��Kn���߬�]s������aK��m�O^��y����۾�ѱ��S�s�_��	�Wֹ@ ����\�5.0
�"ֹ@`�z
S3�c��c�e�I�8��ªHc�/x��n�V�ɰ��:��d,�"��?�� 4�6<��4�0}��B�ȫ]д�g�c�:K���i�g�����k�H��i�iȁ���q� �#2/�a�L������GI�Đk,4���r9mB�)���I���&��W�=�ɝ�3��-��	]���Vz(�ymgG��<?��W圶�X	qSl��u_��}�02S���H�E{�(��7�_���e^�������7�T���.�1�/��i��Ѵ��u���e�፼��+�$�!iW�ޅ
���YI�cg����/'�E@��
�0��~���N�̃!e���}_�6�C<]���W�ӣ��$�u�h*4{oHOm��*����� k6�{?�>i��2��K]��k9;+�Y^�&����d`#q�w��-����[ J�in[��~���SgJA�~@�����xQW0ʰڬ�&$Ku�M��t���y��/�`˜?���D��{��<g��.������ڠp�i-"�@U#��M�u������
�5p�]���Խ�������TO�[al�����,�ӂgF�@��\a����_��X&��>�m�$�y�:�7yGEA��R����D���Ā�LG�cpq���9v�S�'��E1N�c���{z	?M��wF�u�� e�IW�%�h�0�1a(�F?)yJ�@n���dwU�O�	�MV��X�Ӵ�,�,�U��Q��R�I���V,o��g-��6��P	c�~��f�p�����Q���]��'�U�hڄ�+�X�=�<��3��t �2MVde�Mږ��0�o������������2��`��u}�ۼ�����dzm��F�69�F�؟P���.���\O��9���qvI��&ͩ��<�ʋz�(aj�@�1)�6��S��؂��}���Pn�9�_D>3��FR���E�[%����F<��??�}��t��.�x�#�~<�� l �������,�<Mv��P��ad|uOjKcb�b��,y��}� m6�t��0֍]�ܙ��Z\�(Y�6�Y<�7;�O���#-�0Eo���;��s��G�lU�phk7W���ݻ5B�R8���+C��S��81���V�֥�6��CP���+4��*+���NƓ7� �WI��������mY�H|tԝ��9����X���9�����"�!�W��+����4߽ɵ��x,O�ET-r�ѻ\�M�.��M3T��-�11Pc��U�0r��p�Fz��t�<d�W�T�ēo蠛��)B$�����g]%����B�hS]�U�����'cL��0v5�+f�՞�ǜ�ˋ�T֒9�ʋ��K��IcFnUU�'bB���߇Z�����y~R��K�P�����g��h�p�vs1�z�o	iOT��[��d��aÞ�3��_X��VŔT1p��"鸀�<}��*~�PKBeC�  R
  PK  ў,J               202.vec��a��g�=z��V/��X5�7:щN�Kt�N���jt�K���Nx]2��{3sg>L&"�G��Q�"�ߩI-jS'eQ׮�s}АF4�	�4�i��iAKZњ6��ֻ�ٵw�@G:љ.t�����z8����C_�џ�1�AfC�pF0�Q�fc)g\��x��D&1�)Le�mf�Lf1�9�e�Y�������,a)�X�
V��լa-�X��oЍlbs![t+������.v
�G�����`��!���=�1�s��)��4g8�9�s��\���W��*׸�nr����.�����6O�)��x�/x�+^�&�x���=�H5��l��o��E)�E���������PK��ѡ^  �  PK  ў,J               203.p��y<����ƈa�[L({���S�*�!���$br���=��&4G��$c?uR$�7�O8�;z����:������}=���<����"�V6V   ��o��������$Z)(��Fc�q2XiFV񈲬����;�������S60��2:�����$  �DJ
	Ij�a����>P� S���(�2�N�K ��������" ���
��F��(
&*�i�'Fr�����2�����v}���A��%��*)������70��$Z�������YG�s�^?z�\�	�)"2�FB�ͤdJf���ܼ�;Ŵ�Ҳ��{��=�o`4>jz��l�����y��`�54<�~�abr�3=3����������. �+�+���B!P��� ��i򉚑�n�b�Zq�h�"z����݂�{PBBQ�}pq�ٷ�]������ 	�A&�B�8�&������-I�ÒH�+�v�QY��A�[�*I����_���B�5�[��� �=���UXB�ʃ�@�yn�36Ve�D�@<��������:���F��K�Ϙz�R#��a�"��8��[鬒�wOvl��6Y�����i�cdu�Il���Z�2-�	�P�� ̾�7����+�|�״��<���^��$�.~�������p�,]d��_�u�ڋ�+Λ�	1ا�"C�h�qO��f���`'Z�).]C؅�cO�����5��(���hN����-��؎�r������ǲx31�vS8A=S��DGO���Hp��8: �	Hwx��d�K�_�����Q��:K��0V.�*��a��R�״����#��+�􎪥L��}���yr墂�$���x}�+a��6O�pf���K̉��h���9�Ny��	M��ň�T�Wk�o���Q�cX�%49��6�q{�X�g�msI��C�#H�I���7�������'���m�ઋ
��)�?��{}Ri�UĶkx��*�Q(�2�b
�� ��/Mز�'��qA��Yr,�rPh������X9�T;:�)O�'Q�q6�G. ]o�zu��mz�-w��^�ÚG�hL����>|Õ��	"?���{]o� �^�5��m0�@���#�{��k_�n���"��k��_�Y����cZ�@��Pv��ٚ��J����Ɔ7"]��V1��C3Z��t��}����p�#�
V;�.�W�bo=0J'�O�ֆ/��eY�о˰�q��OaHͷ���j糈M��fB�6j�q�� �7�$���b7���I�)�l)�z{���B�[u���`?"&{��R�8��"���)X��,a�,W�<)��U�f-�,�����*�7�{�'�&dm���4jm�����{�>۴��Zñ|���.�.��L7G2�E��X��r�y7��d0wD	'p���<��44-f�`褜�U�h��5�h��Ў��U%�c�i3gu�K]E�нĐ��R��g�P%��&N��e�yyn�(b���l�������[t�^���Kz��^�)�(�9��U��(������6��\�T���Y}N����-*�xn���	��P�)d��̍(y�������%߷0{[?k��'����B��}���v�j����C��id�_��F�5HB7�"�ɺĎ�p8�_m����AX4���{�urU����~��ed�N\�
v64�m�=g;��yqc�TjS�)g�S���<h�,��p�벉Fi�e�ۿ
��0�C�Mv��_å=77�me��Vjf�O�C٨����m9�H,3�$�ќ�b��_������~K_Ly��ۚp��PK�ߴ�S   
  PK  ў,J               203.vec҇�Na����x_{g�Wٲ�&�l�V���&�l��&���QO�{�t��ܝ�u:��J#�
T���w*R��T�)��Us�NjR��ԡ.�l�k҈�4�)�h�#ZصtnEk�Жv��s1:�uv�BW�ѝ����C_�џd�S!��P�1��d��9cu��D&1�)LM)��tf0�Y�fs���b�.`!�X�����t9+X�*V����c=�XL�I7���lc;;�Y,�.�������� �l��r��ȥqROq�3����E�Kz�+\�׹�Mn���;�����>x�#�<ѧ<+I�\_�W��M��V��|�S*�����6��s|/��#r��W�,~�O�8���PK#V�a  �  PK  ў,J               204.p��y<�}�s�c�4�!W��5r�Ќ�´���ǹ�	�<r䚝HE��(���C��,��R2�ѓ#I��R�����gv��|���_������!�@Ή�H P �� � 	$D"$@����B)ʠ��QJ�
��e5U�2�[k�����x<񀎾!���Hm���)�r�~#�� III�4
'#�#�����s�Z �� p� �h�j�<�_�G@�08	JHJI���P��8\\�������$���U$'fKh�V�b��-h��e&IJawᔔ���%���053�;D��;8:�����q����N�9�|)%5-=�u�����7��9%wq�+j~��{P����������Iwϫ~�O�C���ɩ���f��..-��~������A���-����08���Fm5@��$���	U� 'J(�fW�Jj�?���e�Ia��Ƶ��~1��Ē�/����k@� �̓�k`��ȹ�P��-�N���?�8��G?]nUq��K_{�v��!��=[()�`�ɨS�M^� �ʫ��r���;�(��o�%E?��=��Dե$��0P:�4�m]*�Ў%!�TG=p�(�b�$ߧt���Z�����.�����ì9�>e�LO�	�r&���7�!Ꚛ�/0��4Q��Q?Y�z��?&T�KT����͛>w�����
��LҳЕ�������:�%�(8~=\��趭�Ht��s�z=��l�C�	=�]�B���FM*�ɴ��:��!�����R�/�XpX��U�̯*to��((@���~��C�G���`�y�\Zf�5��
]�m�������a�&9,`;>
ݸߌ}�����UO	�6�h\�)p�`���"�c�?�:��?�������0K�p��s�"�F���[�i���)���9t�)F�?�t@�����M���G|XEʺr�� -��尤�����0Qi�n���k�-�l�4_��9�ʷ|�mgr]���%j�z7C��k�3߹?�*�y���	�4]UB��A���'��.��f��<\+T�pq�?�1��}������/�b����yE���+�W 'S��]��)�x������8;������vu�Fd/�.���z���5J�d>V������i��Wx�����k�<�<�a�c�̕�I]k�/W6�G�=�Oп^�?�a�\W�Q�_��Z�^�zwqP_�7>�^��!�q��6�y�c��.=�<�;r4C�Q���We�����+Ƃ�M�3-Zn��"�\$�}msR�ٚ����n�v�=Xê���o�RH����f;����lv�O����2^$ll��}P�Kj����)�.bj$62]6-�*-�*�BOe�Y�zTU��w堅է"���/��@^�v���"��)�a����'K��x�!X�|�
O�k�!���[*�r99��~ȹe�4r6>%l�+�N�p��5N�̂��{�$�Y�Rם�ip�C=|N灼�c���Qu� l�ݞh��P����Es����$�}�]:@�y��k�7�)]�������I��h���e���2��L#�f�����K��?���()"�Jg	�7��5l\[3@��&�T4Ւ�6����&�L|��_�g�D�ԝ^L�$y�M����bo`dtV��"ϋhr�x���~]�)d�*�����N�]�����ڠ��46��Z����C�kw�]U]�"���-j�in* �^?�rX����#�=��3s"'1e��Nn�u�jl>�U��u�N�M��v3��g��қ-&oD�Cn�1��.X�꫚
3*֓��HSGB���7T/+�������ڋ� �c�t}���ps��� �ο<J'���% �� �x��ClX-�rf��"�PKR�J�  F
  PK  ў,J               204.vec҇�Oa���s���;��[��e�M6ٔ�le�M6�W6�dS�?���N��O�O���D��H�J)��N%*S��9E5���5�I-jS��ԣ�MmH#SN�Ҍ�9G��έhM�Ҏ�t�c.F'�L�ҍ���'��M�ҏ�` �R��:��c8#�(F���c�x&0�ILfJ���Ә�f2���an��t>X�"���]��X�
V��լa-�Xφb�����la+��Ύb1v�.v�����\�� m�a�p�c�eqBOr�Ӝ�,�<�^�������r��Tp����w��w��}���>�	Oy�s^�W��������=r!>�'>�|���k!Ƿ��)�O��/��9�PK����`  �  PK  ў,J               205.i��g4�_��F���'���]%zbt� j� �F�����%Q#	�NtF�(QQbƘy����7�Žw��{���g��9k�CX ����:� 1 ]/���r220)9�� ��f�����fcd�c�b�ps�sr���yK���SHVXL*%%�W���'~WJ��M�(((���YihX%y8y$����0�� � �[ 1����@��IJ�����HH����T��� 1DL"%%!���^�RF�*���-f�ȴr^��^������FQP�s����_@PHXDJZFVN^A��������������#KG'g���n��^�G���}�&.>=#3+�mNn^iYyE%�������ֶ��Ώ_��� ����gf���6~�7��w~���99=;�{����E������\�\�$$ �\D��0���@�U�O|�nIF�3���4�R��5��b����>��������,�������k	�]� ��ߴ���hZ��<�Q��۰ĽK����s۫��>��@��_G��`\J�o��$��I�vӘ����Z���UM����[�5O,����@��`�5�fK̈5�MN����������A�V}%�1�N;�r�0���u����m�M�C�)��4�հ
F�v��	#/j��~/t# �2q����V����&?�L�eǔ��)����?m~��1z����G���Ͱ[�/e���L ���̨I��@��M?�M{Z���$���;�1��cF�$x�xj�����vE_��� �!Ƥ��`Ҫ�rxi�@��I�r�τV����n�D_�t�\�٫<�O^�?>zz���Ѱ3��-l|��]��L�w�)�m�0v�����}8]+��f��{��	��?w]�Q��x�F�Ru�Az�|v��p%��TI�ǑY����l�)���P���S��E����x�+�J�2o��93�9!.o��jz2�4��l(��C�Dor�"���1.������2����)%���\{1?X>������~�tH�����q�Y�h���C�f���oW��h�d��BV��` S}A�G������Ny0�fHx�@��x^��L<�;�	χ>�)f;�#/گJ��C�.<�6�t*�e܃��l2"[=2|mk�v� �{���쨽����o3�I6@v�s�hĸ$�]��O�*��YJԨ�R8��cw�>����5��=IF��z_��|/���s��oGY�c&ώ��pA�]K�9���2W�CW���j��*c��KS���g/��$�ѴՉ�����r�Nm�.���A;�ͥ�A��Y.��9��ϓ g\���`�XFC$�{��p�@�E>fp�jr��n7�,���N����L�vZ��J$&kq:������G��F��	=kZ�|�z�Z���v?~�z�i
��X��Tzm��:e��s�� �oo���t���Iή�m�Q�B=�������ڭ{���(�~J|�����A �5�~�c��j����UQGĳ` w�D,w�x9xI��[�4Nt}��8]h�2ҊT`�S�f�V�
�0㦦���p�s��I�?I�\ه*(I&ݡ��kJK��z�n;j
bz�V����G���l
���}6�O�XzI�	q�~�[³{n�69zV�q=�$��I^V���q`��*|����d��jY�=`Ü�N"��r�JU:��1�9g�-�����Yj��,n��~Z1���H���(8N!˿�j�lwh����qftmI@�a��	@��RۯM�A�,[����aP�I�)X�JT!��"wl%eu��om@�H�+WB�ve�qe5E&�W�/�37�F%}��rp��8ކ<�h6�{!�<�gM}S�ڏzX&9�A}N-	;���f������M>�� +<���))��N�3�fa՟&I�*��$�3��]��
�e�9�f 6��r�A��g|K`.�qK׬`���e�ްx�r4;���h�D������Y��}��.{�kc������[f�Z�uCp��-V�]?�H�r��-6N��q���q��Tyп���
��(5v~5�q{����ߡ&��H���f���>v�Gl����;����y�o1^��+��?������}�A�Ml�����z�C=SI{�7�����a\.ԪA�W���(V�'�#s*�*C���E�	BJ��Zݢ�yz�z@\]�I bl����,�wMo;8����E>���^t���fS5Z���;Pgx�R򹉻ڙ/���jl�"�v����_���p�r=yꘜ����mC���#�}�DH��{�i���+�v��@��^o���V�IΟO�BN	 �60�bi�3�R,�;�A��[n����h~��=��� �v;m�cA�.X��h�z_�@�6�����A�{�)�)��;��{!=ԯ� 
|V���wkE1�|�;*�.
�!]��Ց7�k��+�&�"[E�1�<����[����~6Pk��r|�F����V�e��LƊ'I��R�7b��9�v�9N3WC�T��<d�Ù������k��J�N�=�hn�	ψ�U�UV+<+��I�F�=�սj�.Ռ+�p�ָ��X֢s� vV����C�{��z�JwMr�%�0����`J &Кy����%�7�IқDigm�B�R�I�/Z,w/� �o���LF?��<W�M�b����y$���Ժ�M��5��g�F׆ڪŮ?��Š3xӷ�kn���������ew��뎂����J�E�1�Vws�#�s!�����a�6ws6���#�׬|N�`����9S%P�&�fE�Y�I�5���A1 �� ��=l�K��F�F�Lu�*�n*Qbp�p�m�0�мOack<�Ta%Һg�P! �M{b�k��P�L���%:҂M�ϔ1��Gl�G�5����d�Y�%$�Ӱ���iz���EX/��2R]�y��7�kD���B'm��b�����G�{'�W��!�ɯ�XT��Ҩr��3��.�'���q��7�O�H�	ô-���1����omK�_AH�vF�,M��hǧf����Gx�@���0Uz��a ��"G,XL�nL��&�/��ڟmGΖH��9[�sy�^|����v*�Un׭�hׯ{i:f&u[�˙�ٶ�`�^�7q���O0����x%���_�ɚ��V�h�֛�����`n7�1G�����6��'�1Ҧl�xiW>��ɇ��$'�thK^a��
���ק&�j� S$��"���|i���+�5n���e?ٕ��Ψ�'��>�=��~A6�����c[�2$���h`�~ +\O�!����aV��7��}f����C�xM����~�u��6�:)8t1���q�Zu��Ό*��5���>�l�V2�Dh��<��d��F��H��O���kSC�MꅐK�ò����1�X�?T�>���,�J�5�.�X����i�]=% �8 ��κ��9y��=�X7�:\�P�r��8z��/������Z��v/�ϔq�a�V��)Sp�b�J�yڣB������Z{a���gLv�ho��4M�d���"ˇ�5M�^Vu�D��mX�Z*>0Z�ꟾL�����.��4s��^����N�@Z*}Ҥ#����0��l޷��Ki�Ѫ����;r���D�.�<�'c�QM�����	�凋l�#s��RW{�<����b������>bD����:t��E��e�ߚ��Ev�*�n�_eb���P� UZ��Ǩ�^�X\�ȇ�]�*>V�S^��񯅡����#k�Op�k�J��>�`I�@�ᓢig��No�X�l*ߋ�$rϒM��i����/f{�/��}輞��Z��=ŵ�x��E��{g��4[����F>������%��Q�||C�n�o�ѱ93�H�e��sv=����,m/���kR>M��u�DG���Ǘ����Zd��7�ȡI�w�쟈oib�01n�7S���#�U(,���ZA9n�M�q���q���<{`�H+���(e�Y�Ⱥ6�Z���>��x�Z�.�w�O�K@afX��G�ǫ��8X��>����j��Z�߼*��΃!�rKû¿��r�����9�[�\Ul.�k������۟��l�#�Uہ�+l�V�0,����b����c9NGB��]Eг�=ʞ�wd��'���w.��_l�s��a��f�W�ʤsK�&�_EkO3ʱ(W� |�y����g5�:��bd'��߳���u �0��>������\�=T\�%�ON��*k��~��4�%K�2i�a+�r��Ϥє_i
'�CI��h�&0"~���3�)w�`s�j�BvܐF����Ƴ����m<�2�h�1�Z����\��6�{җ�1����0ˌ�j0YgmF�������#�B��O��OA8ѷ���4t-o���q8]Ml���
ZN��=Yw�/�
|Ғ��X$��to�������J��������		�� �K{���U��;O 4M���z��	�����3�?�xn�h9�-]L ��8
��R��>��k����G3L{Zl5�7���8|�ݜ��nb���r��3�d��`B�<.2��ö~#��3�,���^�b0��k��'���G�ة֑�q�Qے����P&J��.�j�:s��Z�4@w��<�Lct>xX@3�3p���K����7�/:>��%��Q��� X=�����p�?�|+e��]K7�A�����`|�O}��`���]�{<Y&N��e���U��.Δe�=7v[�W�� \���ꌽD��1(Ԋ�.�|�kD�|��7]#����h���`�x�M��=LB��&-�RW�頛FؚD�_���煒���Ւ;�|�g��C�̯A���)��ea�JF/D[�Q�C?����#3�Gu#�9�`�w-�?~�B=oyw&X�o_b����.F�ru��uW�H��ݑ��[s3�W�ӟ1�����)�;i�ȉ<��<�$	m�*�S���k$h=uHw��B���1�8��Z-
�!�#�n��	���Χ�T)ҽ*�}L�&�Ճ�� ;��A����İV9�?��.�������7�B��y�`�E��cc��6n?�͙�s��V7�]0Mוt	g��5Ҟ��99/U�@�v�D���ii����zʟ=�����6,Oy�)��HF[w�(��
�i@�:yg������tt�o�_g��ٳ�JS~�{��a�6��f�ѹ.�{1�����`��R��&�����]a۔z)T% �����hݜ�ͥ�,3<v�ދ��f/R��@�,ji����y��&�l�a�p���+�P%�DS
��"�-3Ȏh��T�����8�n/��V�pA�4�LHN�B�K�R�u�p�؆����p���P�f�[G�h0�U��6�1��Z��Ê�G�U �W����m����R$N�J����ܓf��8wn��݃J��i�>^�����̋ذ�|�2�>]T�D�����'�kD�:�i�Q<~d�y��/��R~��}2��f�f? ��2�_��Ȱx��p�G}Z����=x/L����KV��I��%���*�'rv9L�{ֵD�}�3����b���]k#�1!�N�׸ІP�?��_�/x6?�wa{��'�-���^C���yf^��J0I��}�˝Y�����#��=ǫ����.�Q"씪��ڇ�O-�L�IFC�I	���lWn�hH��oM�R�
|��t��;�8$�#��ۋ��Ҳ^Ye�}�ug�9pҹ�$D�|~*�k��i�B�� |O���U6�;�bg*j)�D�z�J�o�}||��I5�ɩt&���=�7������x!��vx�f�@b� ��-˲�cx����%�`��m|_�J�<����6�0'�͵)�O�Tg����mP��II�ꀎ���`Sd!3=��-��܉>�hc���z�������Ka�b�����<��� I}��+����f#�e�駥iO��D���kx%D�^a�H5�V�W%���b�>qR�a-� �Eco�Q'�¦��N%r�>�X3HOW�6������ݏm�D�g$L�#���E����4��T-�l6�IU��rz'�PD'�r��2�c��г���?��ߜ�����M�	E^̚��QX�	`{_gN�v�~,sn	B~h���3�^�r�����}`w���UR�f3��~h��Ĩ�AYW�C �����H�����ROm���c)�3Tia���Ǖs�&>��UG�W4wtƸ�|��:��oK��o��FMϧ�?H����d��i���Xɝ��q�x)g�Jƛ��+�
̙WBD���p��t�<��}�7W,UM.��B�ʸB����͌�Y���έ�ԕ׃���Wn|oFX�]��� N�4}l�����N���V�;vS��=e� d�$�qn8��v%��  �=����O��tι�l�S7��bR�mVD���·��yԹ>���{���G	��x����@i_Dؐ'�F����0r,}�\��JÝ��>D�ꇴ��Hb%"T�����8��kD��m�,�y2��(���������;����&��+U���G�@��P���B�CJ���8���:�v�EP�F1�Gl�[Y&5�0U#(��'����y�mbꝾq/���N����Ɖ��_�b�����\�&Ri��q}�wE�>�����d(*�V��A&�.J���v��K������n�%C�lX����eLYF�:NG Kwh�W
{�1�Lq~+��n���@1o⇇M����>4_����E���.��(+.tƆ[>��?�\R�z^<!���A<o���r3U$���b��O�i��wz��5	{_@/�����w]��q�9���Gb)�	�/�ΰ\ئ��Em�:�&ZW�Z�P��<���L�d��_�}�3�[(AD�,o���W���[�oq}����b�3��k �`�M\�.�c i�;�z1B���Y%;���q���RA�<���z��*��k��Lӿ{�Ҁ��<����k�T ����4_��T};���;�Yy�8�w��R���!:��D>2�FNN 
������b��/�~S�Et���z�줅�ܶ�#���c� ��=W}9N�/M  �,W>���ɔmH��Cىaq����ʉ9G�޳tn�!�_���;'5�z����B�9Q�B����'��ә�{����<���ʚ`�!�	���a��O~��v��-���ĉ!��SF����u # ����B�v�uq� �@i79�c:�O�c�VmΒq�?�* ��K~�9�k#-A���??��c�OjO�^P~E����g�	�&z�0�q����L�#j���j�EG��U�h��<���v���,�p���><i|�����{�WN$,��8W=���wuVs/h�r��ܚ�𓖛f��+	g�E��_ G��^�hX
��{���Q
�F�j������1���,D�TF��PO渙�-ϡZ��ժ����Ioa'��-_��*+�#-f#֋1�� 6-�M+ �8M�t�`����J�ꀔC��]TSD��x�WH�. �"�L�}����Hr�AY{mIH���@�%���{���e2-���CN�iw�/�2������%
-�r
�r�&�l�l�^=-�4^�A $�h߼$�9[��1m���?���{�j� DMk��cD�ƃ%7F\�z�|�o"�I���f�i�u^FS;Ĩv����^���P9�'��f�`�˔���{y�v��С%��2f,U5��T�^t���o3�FZKPIxj��aEF� �t}��嵳	��)�l��V �`�}W9a�? PK���  �  PK  ў,J               206.p��{8�iǟg��<L��0�r�!�֡!�P/F�D�Ų�	�1)a��Ʉ�"�L�DRD2�F��JN-��y�^��w��k���뾯�?���\��O8�8���  E d �@ p�D�QbXI	qq	Y9i������"�ߢ��W�Q����:z����*Z�&$s]C��G@4-!.!/))ORũ��t	� 
�	\��j B1��P��V���@ap�-��  
�A�pL4��0\VU�!G�G�ѱ���<��M���]�[���b7�+(jhj��n72615#�Rv�wp�����˛x�P��#Gÿ����!:&�t♳�$vZ�O�2��/s��޸y����^eUuMmݣ��OZZ��=�~������dt�����������_�����z� �O�_/���Aa�U/�� ���#d��H��)��I�+{�V7p���%�q��;��U�����X�_2������	((jX�u�E8����`��֨[S������!{�h��7��`@�6ˌ��K��t��^u�m������M���1S����/��S؄"*����-���j���P��Z?bI�z�e4��G{�������@?E#@�A&��k;S��s��(ᶩ����/�5��������-�N��$H5E�<��^\6�@ಁ�cz{M�q���uT�@SPJwMo��M<:_��yL�`7�zm�p{`�B��َ!o�q��B ����K&A��3��8�y�Pi�揕��_
�CY��h1�b������Q��XJ��8��Z�,b��[�Ӟ��d/�<��_|�X�?q'*���'�nh��J�� ����+��p j �\h휡C]iGq|�,0R��yj�Z\=�{���l&.%��J�,�lj�]����t���K\'JJAI3!o'��X��+�>��p	�Gg��oo���v���)p�<�/��]�͵���T�=*�jM��� ������r�L� Ǘy>�x�q:��3������u�a| Z'}�6��H?H,W���	��Gl�5�H�hy}�e�l7�䡯cd��ÓE/u�'rv��e Wxz'���F��d&��Ge��2! �|q�A�l$ߕ̭Ѭ���)���(5��j,��E��<��rә�yo���W.�]����:��a�:����7D�u5��9.��ó�guo��mac��q�w�F�=��;�8w�/��Mr-J��I��C��y9�m��:,��[!���j�~)L��$��r%C��*s��c���^���?GN�|ι��f^��@k���s?c��tL��h=覩u"摒����KVS��~n��헒�L������qWF�J4L.v�y|P�cܺⰸ��Z$ǡá4d\�<���ʙ]QJ�z:��SHκ�����?/Nw7|-h7�y�MQ11��ZX �Ț97�O�Joʝ�X�p��!�gR�kO�Q�N���D��k�I�B�e�S�Z�kfd���G5��zn��.��kP{?�@�j��Q��WGF���,�Y���Ȃ���̆�Q���{sr�˷O�r�U�N	V�������+&�
�r����:���Vu^�mVg'��l�a}�;3�6a~
cv6�w�3p���ޥ�|.��T�z��L��Y������Z#��{���J�*ee��CQ��=��VĜq9$Ր���ND]C S�ߩ�`YtC�u�G%��O�溷��l���X�K�Y�g�\��n�Ν��A��Ii�i�D�7�^'���.E!zg�7w5'X��
2�,�,я*�4?g�~ȯ��,�Q8<�Ĕ�x��qdN�8-$C"ۂ|:Tiza:%zI��'ʃDӒ�`,UK3`�5���s�n%FUY��A��0���l~�M�����Y��ҧo��]N�T\�^��c�i��f���w�5��^&�-���6�ٝ��6� ُ��9�,b��{T��q_��������mt�J��-��R�߃)|�/PKS�T�  �
  PK  ў,J               206.vec���Oq�������"{_�le˦k�&����l��&�l�ɦl���=ߝ^�_NDV��@J���*ըN��EM�Z��ԡ.eԣ>hh�Hӄ�4�9-hI�T��vm�m)���@G:љ.t���AOzћ>����@18+��0�3���b46ct,��&2��LɊ1U�1��d���\�y:�,d�Y�R����d�Y�Zֱ�y16�&6�ş٪��Ύ<������a/�Ri�����!=��r��6'�$�8��r��\�������r�����-�͝Bw��y�C�B<�'<��y�K^�:�x�oy�{>��7?�g��|�L�$��B���g��W���Oe�PKu�S�\  �  PK  ў,J               207.p��gT�Y��i$� �"-H	��ŀ�tDETt�:JCA8*3H�8�DA�#*`� ��(E��l���~Ydwϼ�<��=ｿ�<���H��.�.   �$��3������p8�DȢ0�(99�������	�����35��3������b�����R�����`ojaIXmB"�(9����AWK��?��@#@;�� F� h��1�-}'���?�@a2pRVNz�" A `(�B���� S�5'�(�����0��97�N�G*^S8�����F5u�͆�-F�ۭvX��:�"����{xS����:|��ɈȨ�cb���S.���s�~��_p���QRz��6������n�^}C��斧�m�/^����y-ML��~��_X\Z^�п�?r��\`(��r��ѫ�P�����?��G���8��d?B�[xM���wȪ�,�WѾ��w`	��_`�� (Hj8SxF6C��whce��! ���F��n�L�ބ�X�g�Sؒr{��3�r	��Sa}���ۣ��i��s{Nz5h�W`������<��Y���0Ǣ�mRi�mA�[T��a�p �j
3��S��#�����E~5�!�)��!sK��^�f�{{&�O�Dɺy[�6X�	�L$�0{Ak~�E�=�����}��Ͻ�Qy�o���-FM�س����#?	���tI�2����wd����!���[�}���5�Vy$,�j�ٌ6|�gm�i�ͼ�1bJ�N��ӡ��t�/�dXC���}X�AnM�]v��ω�S"f9]�*�C��V�ڜ#��א���Wl�����Uf~�&a����޽1�m��+��C�����"��f��[�r�r�N���s=��="���vy1�ɠ�L^'M��i�3vɳ#J_D�h��80����I{�r�a�}�R��}�<,�e�SI�.�����w�TH�KM"���]B7Ǩ_���B��c�� ų]�ʤ��G�� z���?=	�6��͉�����ߥ����_�w�+���'^B*����YU�Vw!^��������Ɇs��6�%�����n��(#ҍ�xu��D~ޓ5�g7�7:��1��,�G�d�Tw^��8�w������2�z\DY��j�0�x<����i�����
K�k�~�ԏ����`���9�h���VDoO��d����K�XH�<�]�i3W���n�2f������+K^\6Hb��lQ�,�է��W�2��@�� �!�8a̓����³ͦ�h�����Yu���[�}�J�����<����;��?�X^�`ݻ�T����Ӭ'5��g���i�'�CU'����|�^m��
b�<H.��#���F���8��c����u��J5��{����qa��z��F�5�a��ѽ�5��W>/`Z��xk1�;�4�4,yr
�@��"�n+�g���+�ŷBwt���PK��J�Z�f��I��Y�>Qf;��q^�r�[������)�15���7΁��ޭؿ�xr�}u��`d��$@�K}?�aV�S��t;�FL,�Go[���3�7֛�eXG�����-�:�j�N\����y�K:/J��WZD�H�K�A���Q���v�|�� �z�^��$_=͍��%��b�������:�[9Y���&O����I\^���j8�}�{��;�jX3T�u�Y�kE|5b���s��h�.ݍh�=D�U��o�јĥ��[���c'h�� �EE���e�{���������zD�8���s�t-vϒ��N�< kk�g����j���7'�>��R'��M�F���L;�h����_O'f]N����u��R���c�%�H�9a[�˹P������8�bl�+.����E��LS�_�� ���-F�{��+O�������31'k�$ ���\��ְ��50\�e���}N�g����Zܷ���?PK��� �  �
  PK  ў,J               207.vec҇�Na���y<����.[ٲ�&�l�V���&�l��&���Q�y�ۥ������t:���,2W�J��2U�J��Eu��5�Em�P�zԧ�MCmDc�Дf4�-S)ZٵvnC[�ўt���BW�ѝ����C_�џd��Bѡc8#�(F3�f��c<��$&3��Y�t:3��,f3�����c�.`!�X�����`%�X�����t=ؘ�b�nf[��vv�3�c��f{���T�z�C�<��r��HeqROq�3����E�Kz�+\�׹�]o�-��z���<��}�G<��<ѧ<s~�/x�+^�&�x��x�>��3?���|�H��G!��H�+K�;����oE�?PK�=(F`  �  PK  ў,J               208.p��y<�{���1���5"32�#7�jb���ZT��I�ȸ)&#u͍,Y��qu��C�2��[YF�%ۨLa��׳��\�����>���~����=����a��^  �� �~�@IH %($))�BK�2�RRҪ�
r����&5uu-�����!V]����vcSSSM]s��&�FS���@$%%���UddTL6�o6��M� `P��@�@1"j4�y" ���A�08B��DK��6 P��8\��8!�٘(�@�Fj�MbS�Q�=半��s80�$ZIYEUMg�.^O�t��w;�-llI{���;�p��<x谏�ɿ��;�~6��㹨�K���@OM�����u#�q�nAὢ�_*VV=��a��M�O[Z��;^�z���ܞ޾��軱q�����`���OK��_�  �/��\1���_� �ȯ8b���<���>��m����7Jb	�s�'º�J8�a���h�����"�7��� iD�<��XxF2$��+��@��T�5�keJ<u*���ګ�ؕM
̜�F��:LHWF�_����a�N��zq3�$�`���`y\ɻ�J۠�_��.u\��m>e�s,��ae�?�=���X���,���+�v�-k)p�9e�cq#2%o��|r����L�\1/��N�E>T�<%�$�$��Bz���B�U��v-�k8ڛ�R���kQ3u�ӠE�S#� �Y��t��"�z0�W[3��/G����d��|?��Y;͸5%Y�ӧ�����B<�z��cF��?Oek���5��Z��2u�x329�d|�wY�<O}<xx�J��Z��I"h�%_�6��`w�~�����(1$�w�d��(++u}�v�9��9�H�M�+#��[X7��ҁ_2D���h���n���K	Ez~�:C�q<aZ�+�����1����u�~�(�aVϤdK\ޛ��"���kn��[���/=�B&������Ck~�{�O#��
�C\��D@��m��9N���������(�Լ�� ��X/፫z���O}�̊F�ٱ^%Ѽ���n��Y���B����b'��`4�����u����O��N��s��>����sX �e�-X�Fzs�t;Q�55���_v�ȹ�]�����ϗwz���ykuݭ9SY�_�S =�x�X�=�����Z�yV<��S�	{z�r�
�i�T�6����v��j��ʙ�T���FmF���Qe�]���+q�m���>�3�t4�qq-Y�q?�U֌�7ò�����e������5y��nǝ��r�U�W��3l�ۚ)����3��Zz_5�c�JRiM�x�%jeڇ�D0V�
�x�)�����Ƥ�Эߺ�nz>��ʄ-j ���{���x�1p��ұ�|������ ��Ap��]z��(�\�o
O�al��woԝs��R�����Ś�z+mc��n����d���������WP0�����#~d{�Aڐ�]\�a!�p��[뜍�a�D� ������#ۡg��bU8����sY�dy�e�m!�cp����^�Mz˛�;v;k�?D��K�;�D�8�x(wqB�qp���]x{�ڰ������v �7��5�q]������7
�E�|�A���>j��+_˕h��)|KY�칶�N'3�3ev��c|�܍wJ����c�Q��W/���K�R�Ĕ8����#Xr�mKg6�g�c�����>�"����k�����b���Τa{oް�Ȇ��i�
�W'�>	�jٞ�~���Ӟ<)~��z�4����s�f��"�Ϥ�{x����*�VŢ�F�^��/�

�}�W�jjgc�'FXIl���V�ϊ�^���@\H~2�6V �0<'�*�bçb\����_�8iַ���Hz?���{���>O�S���v�ug��V�I~vk-@Q�? PK���  ^
  PK  ў,J               208.vecч�Nq���y���޻le˦k�&���M6�d�M6�dS�?�x��K�W�_�O��9YYd�%���N%*S�����;נ&��M�R��6�!�hL�Ҍ�H��]+�ִ�-�hO:҉�t�+��Nzҋ���/��� 2(+�`�P�1��d�Y�uc�x&0�IL���S��tf0�Y�fNV��:��,`!�X��.ѥ,c9+X�*V����c}����&6�����6��������a/�RY��,�qHs����	=�)Ns��������E��e�p�k\�7mn�m�dy��{��y�"�����%�x�R�ѷ��=�號�3_l�V��V��{I���g��W����?PK���`  �  PK  ў,J               209.p��y8�����a�2�H�b��X�c)�ʱos�0�B8����i��hl�5�yD�H4���X�VSq5w���{��G���|���}�������wm`mP�k�d��  �|��0` ���R0��FȠ0�($�YQI�EUSc����VmCݭ8-uu�����1�H��%��	V�����$ iii�"+�Bئ���?��c � Y� �A4h�Д�	��C�0)8BZ)�P� �A
���P��i�: E���H)��8���}����	��i�
�I��Qޤ�Yu��.^o���̜dakG�wpt��~�����a����0��G�c��	�O��t6=#��J��ܼ��]��-(,*.�s�^����yu��OZZ�ڟvt��|��/NLNMϼ������ߗ���׽@ ����^h�
�@��^ p��4��XJцd(�)̞��UM�Z��Dؠ���6qt��u����;�����_b��P��� h������0���@y$�m��z���_0L,E �N>��
>�>�;��b�B�8Uk3�`9�Bs��3����+�K���l�;�~+����|�CYV�[�O;�O������g�D.�O`��kM�9���dQv��Ȟ�x����h�0t���ƴ��q�ZҲ{��Faט��sY��1��|L����y\`"$�}�\���b�ז˭reZ,"L��q����SQ�ڙn��b4ut/��k B(����ɗf|�]#�����K�>�z3�Ǡ\֎<�̟aIQ����r�����(��"��{�9]�*������%*$�����%:̫��,����Xk�
lD���zœ��/*Q�S��Uf������?0�C7!�Z�I3s޼���(���Ih�1I����l�r��~�|e~ ^�ؤ?����X}����3�ӿz���� [Y%��^������u�R���Q3ֱ��ާT��&�iY�d�s�X\����)bj�O}�:u��B
��,��q�Ϝ�ӗw��B~/������v�}OFc�+�t1^���zƢ���EޏҪ{3�s��`#c![�(���|_�XCW>�������ݾ}��֡t��=I=�~� ���~����3Rw"��\���Ш���@v'Zz��8k�V+]������|����/w{��ZР�R+IPzڲ��1y���OD'\DX��jF[ӥ�a�;4v�|�#6�����6�4��6ww��y.�@*��p���`~nB^n�ы-�9âr�b�tOਪ~c~��@N����^^�i��̣:��,�
��6 ��KJh��{}�k��+q�_|��Bu���0������c���E;�6�
}��i`��+�7�hh�Y@�)�K��D(�n>]�:5\�[Wa�󽲳J(�z�v��7��LiV@�7v¢����!�Io���M��:�����N7(��Q��W����I�I��購�-]���`{��І�"a��ս���Rɐ�Iz�U�8�zL��7bw�騩�Ѩ4���Ζ�f��om��f'��ծ�����*��������h9kH��y�t�Qo�9,��i�	����~�G՛u�=�Bc��oy$���"2���Dr�%]6 <�r�~�ԈQV-���`�rk�1�N��U���Ց�~ƍ����,�:��nqv�$�(�]����"gc2):�U����>��Яy�Z�,/���d�_1�y�=W��l��8����V�M6�*|+V�(���e��PKޭ��{O�S1�}�L��~+d4y"�(��>[~yh��N��	��vl�4�֌<�O0#�1q��8Ò���赩L��H(�r��i�!O���*�g�	��X���)�B���pT�2�z&�>�'}t���y�p?�Q�ue{70i7����[Ŧy���X�[q�B���PK��ë�  Q
  PK  ў,J               209.vec���Oq�����{흽w�ʖMזM6e+�l��&�l�ɦl�q��=?�^?|:'"+��S��R���De�P5��]u�Ԥ��C]�Qߦ�6��iBS�ќ�o��k�ܚ6����@G:љ.t���AOzћ>����@e��C�0�3�����f��a,��&2��YSt*Ә�f2�W��s���������,a)�X�
V��լa-�X��A7���la��M���f��b7{�c��Ke�_p���!=��r��6'�$�8��r��\�������r�����-���r��<�!�R�c}�Ӽ��9/x�+�~�R�q~�;��Y��3_l�S|+M�$ŏH�3K�+����O��PKruϓc  �  PK  ў,J               210.i��g4������A2�F�6j0�"z��hѣG��'z"H�����.z�Ę���nys_�{�������{�}��f�f������� ��n�� 	1!	111))	��|����%��������1;##��� �rIH�I=���<RRR�0��"���*����V��O���Tx *��N z�NB���?��" $"&!%�s�P{����	@���Q��8@@EH�*(GtO�-1�3�P`�7v��6Z�a3� R2��z·\�<�pQ1q	ɧ
�J�*�j:�z�/��-,��Y�غ��{|���	��D&$&%�|NMK�����_PXT\U]S[W������������|brjzfvn~um}csk{gw���/������?\x ����Eu˅O@ " ����$P�
Q�i�u��&HB#�����]X����e�����y���&����"�_`��k ��n����}�O-�@$��*y���j�	m�1�h�!�O��݂�*x���X�����v� � ��G\s�j�p��=�{�I< zα0����!ȩ���n���Ǻ�����6Y��F�GU6Z]-�UM��ͯp�a=|�e&�Q��U\�2�K��ѹ����Ӽ6J a�xG�q��б���3OQ��y#���rW�F۫t����Ç���c���	Γ=nܝ�'�uu��
|^҂1v���ʴM���u?�>lgq��0�ʞe�>�� �u�)�b�����WџwJ}67��������S��ԱOAo6�{*�N�ea�S�D��=|-z�����Iy^�������ɡ��x����]�E{d�\�* �����g��݁�2�X��*�����M�NA|�Ɇ/>G0�1������3-eׄ��<�]��H����>�7 Y%#���9��(2XZ�P}����w�@��dʶ����<
�A��vL����qw{g�U��f��yZ�Ժ�,	-X"*�x���?�x:�I��@�UN�K�̜*.ɍ��v���t��ݺz����Ǚ�2a}u�N��G�(�T����EWȕ�Q����T��C�oDi��=]3�۩��?v�sn������̝�o%<���^�6n���Y���}���XY袶��ߐ�"DŦ���w�~���"���Hq��I$�+�>ϸ$�pn�����+�Tf�P�	�݈�f�Z�Ɂ�(A<�Hk��ad���U�/c�rv����()?�(���U�,�-1^��Į,�)�m���p� ��BY��/��j�d_��m"��~埙��/��)���^GOj��k�z,�(�x�^�������K8����k��M���D��UY��u��<|B>H��>�vض�/h���V����jD9��E����v��D�����Rq��I�>"���y8	���z����I@�NZ��s�ɔ�6��OR�������������Au�+�=�X������앍o7���-�x�2�L�~��iG|��'R�+���TO�S3�T���=��؃0е�i�[��+I|�{'����
��U�� ,�p]��,0,�5:�0��������ۑ	t:H��Go���@f�/i���ɮ�
���f�o�S�Z��T�b�ь�va<ٍKMC�X�
.9��#��%LZ^��#bj���"����(C��F�f�s%�-�Y0^\t��4��W�އ��L��5ۭ&x�F�c��¦�a/?E��,�@e��B�H{þU���cQ��������Z+�WI�.Y9\r�#�$|Ue�d��R���d�ĉ�ڟ��/��X8�~�p�C�q=��&�����!���R���P��L��|������˵���?:������!��`ݩ5U�j�0���,Xח�Cn��Ec�'���U���[��(^��^r+J��R7 �4��k�NE�d�ߚ��ۑ�FYC`�Q2u�׭�!Lg�~Yy��G�0��H-��؁GX}.v�#0f��U���_���/��OZ ��[�n V#��O�K�Wɐ��P������8�{G]�m��O�s� qZ@�$Xk�>��`'&`�u�u={�1@�F	����O�Hl�GfN�m�!fN��E���������ͪ�2�.�"��[�O��Yn*_��8R�������(�҆���?�9U���I��n?~�����DdR��Cy���|��֥�R�KE���]t�����i�)-��Lr�ч_��^��B���d�+�Be3��p6ߪqǐe_���^x�A;���f͋f:JU��G;����&��NǦ�4�.dK@��c`ɭDM�,�{#��ƈZ_�;1� j�	�,�*��c���i��?V��YC\~�t�9�%w5�wzS�F1/����ɀA������_8��\��Q|H�����aK�=�=�C�Y:6��D���}6�mr�3���q::�v��e��]��;[��=p!m��\��_�l�#�8tj9��W#G�Gֱ6''��.�^!�AXr�J��wZ�4t�����ߍ�{�{�Ct��JM
h���d�[��s�]T�4��{�]�>hJ!���	����ȹ��#M�Ub��m#C����:mH��Oh�m"&�Sf�y_��*�0�Or�G�!=�Z#8��D�h�<�L��b���^=����Gy��aM�:�n�F�J�66����"p��x�,�&ۆ�G?�ShS���d��Օ������8��ou�X�M��g�Q�,:Q���˙��ϗ�%l��:����4_}.�����!��~_���ӓ���RL�{zϐk�I�y���c��	��W�9٭�#gy�=���,�6-)
W�4O���E
o�MD7JB��Wz*��Bz��ˤ��J#i=JB�$Z�6PNꇸ����2�����Ow�t��܁:�_!�X�	����sJ�1<u�G��ǟ�wRz�9\Yc�����L����A�h�=:2��)�#!2��Yi��QX�t{��� �����_��v	k5>�8�Gd�-Z
��XF�1"�;�� ��(\������X��e��ޤ"^��|���\t�(J����gh�gէ'׭Q��.pr�(��&�_�6���W�y-o*-�b�@�B�2�=��߹�R�^u�L���=�Ѕ%�X��@�`/�~��}.	�ic��lTQdi�Q�P'�K@�B��#tp��r��zU�=�&|�#�姌�����Hzպ���"���4��N��l�^�)�g�+^v}g����3����W[���7�l�R:���t��ў=^ �tA� ��^���Ib��H�Y;.����y��؍ ��v�rE�e���~�6\���ni����^�3��\A#n *�T���`�W���N����mJ��Մ� 	���y�a�Z��Z�,����r�^N�x�թ`"�_	\�p�d@�ǃ�������&<D���˅0�+)
�G��/�P���?��'�Qy���!>���Z��
��e���R��R�C׆��G�\������b�{߫����f�l���:x�U\�[}]�-�m��H�̊�J�\�d���C)�U�Y�c��ޥ@$RP�ma�ݣ�CP	e{�Ӂ���`?����P+��t���T��l^�,!Dςk,��9�</��Ő!����׃�n��jcyp���aE��H�#���5ˑ�/�̉rn #�GC&�eHxӃ��0=���0�jL��Z̴BCͯ(�ߏ����1X�G2���v�ocW�o�l��S��/��*m�����H��<J�~��D؃��3r�xb^�<}cN����ֱ����}�H>�����m��Җ��?7bwѓ�1�v�b�������IEi��_�{���5�m�)�X�/d��/K(�x&SK�m��~����M�@Q���SG���B���Pz�5��]�m��;���U��ul%9b��Z��v٫�Ύ�=��2��2"u*�I���H{��r0vaw�����FD�or8�Y���-99)���SŚ�R���g.R���+w��}��G�|��}-�H">e�;9��U�/q�����H<�cG>ԘJ�<q��5��t������8G���#$������=߾�*�0E{.�n�<ND^�O�t%�I�k��ʮe5�y�`��K�E�y��=���u��S�#`+� D&ČABz��{�z�_�����	�G�����mϺS�J�]1�/��4��l���<�������P%Ȅ��(��-jCLJ�p䶎4��5��_��+�k3�tҚ�_��F�{�}�ӏ�nkaJL��w0r>��(��1�,SD{���P���͌Ȍ��keA%��(�l��z��β�C%���;?��v�\�����Y���nMYϤܳ9ڰi}���(d��qڷUZ���Q+t��^wp�Y��B�?;��?���:�>�6�j�b�c���i���h�~��e��6	�_j�2]��C�`25"�_*�[�[�ا�d;���J�*RĽ���Ԕ
3d�N�Pv�{Œ�Bw]�ڞ���s E��`�!D*O��gx1�����y����t���.��FOT�W�b�K�:�A��gׁ��!\��j��?��}�f2�ǫVg@_��|O�Ͻ��_&�:l�9�-���gW�S��]V�XH)zrtQy�1`������Xi�`�D�y�S��
� XA������3���^&Y4r}DG���Ó&������m�U�Vcaɓ}!�-���'ϼ���8���z�4�����h*���x��;SMs�����Fg)zo�7S�Ϋ�����M\-]e˵�j0�cF,����b�qlO�(�h:m�uf�K�"�K*� �������Y~7�.��g������c����C����w�s�C�]�ұ��֑�-���ٶN3�$�3�+K�����G��#&�����nl"�\���G�O��$�!}�3��;����p��9k���ڌ�հ�s������d�-�����ڀ�#IһQ��u���޽"�i�'l�o��5�Aç��/H7V��S���R�D���c���%_y-��qG�2y�7�Z���V��6�E���#C���9z&���=�<#g�*e�d��È>�F�z[vu���D�v�G�y��nS���_�^8Hr�q�Ň�.Q�H���O]�@��̇�ߎ��RX���GH��N���|~{4k�棬`Q�=R��E��(=j�$*G#	�@�����;���I0�X�fp���"��y�� �nd���D�[����Q��Ҽ�ru%ip�r�2%��I���W�~�<ь�.Tn��'�`��QV1�7M�[�h�`�6��.}�dhPp���Eۈ�>,1��0i�n'թgt=6��F��}h/�<U���OP���:�G�{W#c���7}v��;Ǖ����h�����퉒��w��H�A-����):3��8��s��oqY)�W+̚���7�4���yꎫ��ˏ�~.[r���!n{pz����/o#�D�_��k?���_�$���9)�;Ӽ�?3Ѝ	��B�T)l[ ��K�r��1���!�ђmϐ9��Q�����ZIL&���M�0}uk2$Z�Ö�DL�.�>s����8�tc+�^��4��ay�39��گ�ӽ��B��߹Y��݉�(�p�@H�����g"�p N"Am�?ӧ�1 �\��91K9�ed��|?@z�����?�S��ǖB<$�C(�oI�ޥ�8�ݸp*r7[�y�ӿ��Ċ5t�0�o'm�s|�$lYZx͜�b���4:'T���T��|ۡs$O�����^�����~��}��ATv×���/��V��ZE�a �?Y�L.\k9	�/�!ڱ��j��v�ѩ۰���wD:���]MB��:�)w�%=<�n�}�*v�Vt�)���×��F(/�ެ�b�D�b�ݸ�9�,W!A(F(�s���?���k��-G��ț�r-�`���l�) Bo�&ՙtT<�]�G#_�xV���grލ.@�sVu>�:vB���?������WсZ�o�2����V�}�9�����W �	z̐.��s2(�j�bk���> �IʠyT��~e�c����nbol�.�k�Cmzy�q>5�q{���ZC6�{��摨��SX�(,Pa񹧞���h�TK���[�~:�Ⱥ���͡ _����X�ӛA������䯦沝��ȃU�_H� �h�f�}���}7��-C�#�!U�H�.��Ja�i�/�v�d�g�7�|�f���O��k��r��a^(. ��;)��ůKb+�o,�k�SNg�AbZ�S��7����K/_eEz2c`���תX�Mh�@)|�W�?�f�����_�����`7�8��mpYDld2t;�Ǧ�UP���g2�>0����:�b�9��5�)W[R!;���;8�5Q��@���{ly�Ra�< h ��ũ8=�K7$S�ۆ9�t9��Ɔ����#���=�k��Rȱ$x�$���S�<&�B}}<;��/��؝���FKQ��%�ʟ���#��$��wj��A����,��Tqo�s@d�x���ݔ���O� �6����Ga0�q���6���檺���쭭�Y�Y�Y;�GㆈE�[���p8������ՆI��C�g_ѻ�\����q-ҁ�;\�_f�<9e�;~IIH�2�5��J%�O�=���(��F2u�ˢ��Ft�]��#g]f�1���^q���^+��
f؅�=�%i$�]�Jpe��
3wRG�ę=���n���.��?�Y�	J@�ߑ O���ZH����@�����]���w�5k�2Ф�#��/.҆������P������ۼ����Գ������EK��d�����X�D��:Q6� ���jR�Gs&���h�P������������}PE��<:5q�:��h~`e˻�$�Cr^<��
�K�}��"56����M�8�_���Y��̛U6���e�Ib�G\7@��ض����Ʈe%����LD��HSɫ+��BΨR��D	V_Iv�#��#���3
�X-��BB�#B8~��Z�k��xn�f�f@ꢊd�1���8x�=��q������"k�q�[b=�s
����cy� ����'gb��^m���T�Ƙvن�6�hj�1;u�	�e��$U�uI=�*S����׷���"g ^���wk�=0����<���|�2O<���66�t��V)�=/s��*H������sl��璔T�YbC�ɻ�>��CF�<��&ᅯ����媽��' �X�3�>o&�)L?�E��6W���u*\ɝ�����[V�Z=�v�l8��� �Y&BIcR�;�L_� ���,WLi{�Z�v
�su�U�Xnm@��s���۟S3Ox=�97���뇃[�1��D����:�o1�yO�y$�� p<+�
)Z'>�9�on�Q|S�}�b����m������|�F��g����?
~��i����
�A��`> &�|�0ޅ�t���泱׽3c���SC#�k�/�q�w��1\a8[Xih�Rq�@�nF�)`)��+�4^��D���CDZ��]�C<�1>���nc`�_��4ߞ��$�՚h-~�����@����D
�h-��Lv���@�|ŕe����:$��X�,p�?YU�p�%���úgW�Zu�0���AǳdY�#��u-���8Tj�v����c�d��_Y���&`W�Xk|^m?Y�!N�B<�%��d�xL{���9���PK�zs�  <  PK  ў,J               211.p��}<���{d���F6L�Șې{��S�La��+�"�R򬓆ɭ��Fn�I�t�Z��1$E�V��z����������z]��}}?��%�� \��t  �t�� ���a�222���ZQA^^A]Y�ވ�im�jj�	&�x�ͺ��DK�ͦ$2��ӷ���m51'�};�@ ���̴5���琴(Y�P� `�I���N�{ ��edr��� 0C!0*��H� S�&m��0dt�h���"Y]�����y�y '!��'5u��&}��!��K����v����e��瞽^�>���>�=~"*�lBbҹ�^FfVvNn������\z�FYuͭ������wtv��~��i�������ѱ��WS�3��X\Z��I�������%�C���7.���((L�W�Ɛ	`���ɢ�Ӌ��"t���1��>9UyTo��w��,��"�'ؿ���$mP��F��Ͱ�#��w��i�䞬B����|��
�B�P���ɴ�{�~d��,�`"�h~�eDA^<�X������I���t�&)�F�&�T��[N),}k00�]hh�����e$j�|��k��S/�J�\'f6�R�P�=�"N9���p|���/�,�5ע�5F�ma��G�����Z�+��+�YXu�\�5�u_=dJ.ޫpO��pS�O����qB(S%����հ������61�l#]'�,����=�z�����p}AAѪg��Raxo��MTϠa��ih7��̱1��Q�NBF�2���+�+��y��x�ǐ`�k��0w���.�}�}4��A�WK��? X��ϖ�����g��@e��h��ȸc$��P~W<rТ�P,�zdoqe�-ͭm�.Nu���<�����hh�`T~9l��D�3mN�A���s��)c噿s�C��$'���=rD���d�C��/voީ�DV��E�W�^m�a�>�16	4 ��	 `:�v/	lP߆��.�x<5�7�]1�>�ZGT���o�=A�fd����(�Ud[m��	"Kך�a]�SSgRnh_���UzCҗ��_�|;�*���I��BGv��b���89eښ�j���u�Cܥz��i�q�]u;t�M����h���q�W�_�tLw��L�qͯf�sk(j
^q.�7�؋�xU��rocK�:R�tiۜ<N6�x[ɮ�p�c�����d�uw⼋0W��
��
�;!�/.p-c��q�B���ܢ���]��u��H]h*��5�h-�i��Y�ʏ�Ld�����S�>���P�;0�tfRX�R'��Y�e���'�^�m��Rw�QL1i�d��J�7�	�>��,~}}.�a_~͵j��i�؆��)��˻B�q��T4��z3����>U �����h�XVAI��؜B��sG1�����Hm$
��v�+�=�;�]g�m��aoX��r���}��{Z��U8�Mm�_��Pp	S�����{3����x�ޒ��>L�걡�F����Ƚ���;�v7Nk�D�znqVQ���ˈ��֒��ϱ�[��q�ر<S	@�y��S54�HoU��O���kj��������#W^yx몯�_��UWf�XVl�)�w�q��3�$@H��?��(�XK������i�?��N��wӻfyo��#qrP���R����Rӵ8N1}S%@P/XA+���N�j�Ho3�5�ТJD�$���jB�#���q"X�y���h��қ�1+���i���Q�Ryˣۀ	�N��ƣ�.�#$Q����$����Hϐ��e~��>b�fGR㠧������F�#Wk	��<>Bm]�Oq�#���#0?O�K�K�_Kw��h��ںȄ�K�8��v��Pp�b�/w����g��O6ً��Z�A���Cul�ob.�[�����I���!O�e1h�k���PK���  �
  PK  ў,J               211.vec���Oq����~�w��e+�M6ٔ�le�kg�M6�7�l��G|<tz���=��9}#���\�����*T��S!j��t�Em�P�zԧmic�Дf4�-i�~Gk�6�miG{:БNt�]�FwzГ^��}�GP�@18+��0�3���b4c�,��8�3��Lb2S�j3M�3���b6s��<泀�,b1KX�2�����b5k|�����l��ب������6�����f��b7{�˾T�� S��0G8�1�ۜГ��4g8�9�s��^�2W��5�{�z����g�л��>�L)�bI<�#�8?��y�K�W��7���#���O6�����[������:����PK�:�b  �  PK  ў,J               212.p͔y<���?3f��,#�h�ap����X&�I�ҡe(9)ǒ�Rɚ,3��HaP�vYS��E�,#K�An��8���.��ý���|_�����y}����<ۃ�� !s�c� �  � �o ��a�8�D"�P����"��P2R�2Rh�,N]I�*�F�+�������Q�����S����)"�H~	AA	M9����u�04�! �!��v#�ᾓ����@yap����P.�����roop��0����LԊ
�z�4��3��%�b��8-g�$�~q	I)E%�����C�ut��%��Q��ۜ���w8������~��s՗v��? 4,<�v䝨��Ĥ{ɬvfV���9�y�eO�+*��k^4465������}��?0��x?9�����ť�յ��_��p� �G�[.a.
��w�@�k;	�P^9�����%��F���3J��Z�b���|�q��
�;h���3�����`��  �� � 	X����xQV����Q,���Ir�@�B�ګvS
"b����}���ֺ����т��W
5�\�-D�?�D^���i�Q|�ZN�<?a<�����꘩̭N���t�������8��f���P��9'�:��yN^�AԊ�jFY��?��>���z՞�=B]a��{u���)C��K�]z�C8�b��iwy�)ѳ�&���sD��۷��7��� $�HN�� ���������`bb��FxvTW;
�� e�����`l!n�Uh�3)�P����j�Ѣ�M^�zQb\���]�	�˥�U�裬N�dԉ��0{HZ��U�J^~C��S�J��4̄�頝QJX�����T��0,����U���{��(�M3�óo�&������ġVI("�EQ�|W�y`Iafc�b~x������3]Ȧ���<o>+)2<��g<�E���&vO#\{��<0�f�QS�7�-��.I643�5��2p�%!{�1��
,�,�_�O٧��qY�{��~��U֔�ໜa���o/�}e�Kg�*׆n�d[z�ޚÎ:��\��W�(sz<,M�s�6/mΩd�����si���T�����cV��,_=Ss^�-�>�y	6�^Ęs2͔eZ=H�M��϶wSY��#-u���!�A͵�&jå�w�{���ۜ� �]���F)E�ᥝ��U�A����NUI�j�� S�;�cЩ[屖��+�^�69;W��ȺNX�I{����1��,2�)w�ģv���b�2�%[0b]����i��5�4��ڹJ�x���9�;8���7�h�'7D���ft�<ǖ8�I)��B�;����~��k���ؘߤ>X;�p����O��2tȕ�%�����\�j�}t�2<u"~�葸rJJ>�x{}�X�腦��5��ΤJ,K�a�i��Z�s�G�W��I�:�ٯ��0�@'������zA��6����c�u|H��	n��]��-]e���M�4�EoP;|�`+��?�P�����Ѓ��+"g�EX:�	J���whZז�x4��LMrDr� u�����Z��5$y��*-�l�#!���+!�����M��Vkw?u��%��$H�l�wg���KԵ�"-�2i�����������^.O���>8�d��*�B�Q�ww�Ȏ�8��ݦӬ��>F_����1��s�)�������*C>WhLSZ))�q/��eq\c�������L҈��60v�v7R{����^;�j�q=�Ğ�7'[&�O|٠Ĵ1�KŒo*V�~GC��*������p�������l+���^�M��Q�2,�m_D���VP�h��1�nv88�"y��s�s+�պɛo� +b������Y�/	�Bqu��_l0L�g�g��>*�1=i%�Gn5
;��]�q����>Op�)?!+A�`J��`��iP�f�M$	��b�/��<���PK}�X֢  ^
  PK  ў,J               212.vec҇��q����w��{�͕�l�.��C��V8+�e�M�M6Y��?��}<����ӷW�o}�Fd���rP��wjR���I��kWϹ>hH#ӄ�4�kn�¹%�hM�Ҏ"ڧ?����s':Ӆ�t�;���'��M�ҏ�` ���2���r1RG1�1�e�)aB��D��d�0�iLg3mf�l�0�R�1�,d�Y�R����d��Y�ѵ�c�/�A7����|��������mw�.v��ѽ�c?(O�qPq�#�ǽ焞�9��9�Y�q�\��e��U�q�Tx�M�es[�p�{��y��TO�)�x�^�׼I)��;��T�||��|���7�MUA���G���/����PK�}8!b  �  PK  ў,J               213.p͔y8�k�?�DD{EBQi,Q�v�Xc_j�i/j����4�Tվ6]�����a�ڵ��ZB;(��P��4�-JQ�����ϸf�9����}��=���9�q@���� �  @��$`08L\�#�R�RH����V��������PVݯ��D0�ܯ������ ��L�t�H�I@!���߱C����B��C�
�$@K��b(��� NT�8�[ �P��%�Hу:i@�@Ġqq(Tt-��(q+��8\��ϸ/�f]���k�G��	jBRn�����^�&QO��Јlls��������������S���:G��y%1)9%5�=3�vvNn^~����Ҳ�����ohlj~�������~>�j���o8C�\����4fvn~a�����յM.����˅q�A�(|���|������d�\��/�UI�k���j��eOP�%��z\��M����3�����w�qRP�<
� >6X���Ga�ṵdu&w���ؐI"�A�$��3���ۻ���0�=�0���C*1~q�ң�|z1ģ(�[/;��Q�`�T>�S'��3��{�:;WR��:���D="�U�����r��.E`с�$xb/2mw�}�3=�NUh�*���|~�ο/��c[���{� ��ז{����A�c&�_$�83�Y_mpM�{ח:Ώ8Sc�2��i��g��B�����e�N ��y�9��<����:�^����X�T~R���|ۈ(t�f�O�Kʘvs�&�p�t�í����q>�u�*��F�Y���'�֬f�N���#���Ʃ�J��/���|��ߥ�������Ytb
���#��_�j�K�˶n���2B��y���Qk��]�LV�_'�5օ �6�_��l����vu��m�z��2t��4f$�\�&�?Z��}#���^l�*d�~Y�֜��	?k����U~�v\q�Ff"t�0��P~�Ml2���M�<ys�9r׵��zꨋ��$����(Z�>m"��u�Y�ꃦEy�Ò�˕��C=�Ej��Ⱦ�m����*�'T��e២d�[e���� ���vvY.w���Rw��ԃ���l5�#~CLߍu{˱?P6x�z��ʷ��|n!�z�<�'�][rE�ׯ�3�.�����@�bw:�K���YC�[�S*�r�����)Lۭ��|©u��}��U��O�0�RڢrD�
۶�͂K�ōA��k���4Z��ƒ�S�G���7�	�tF��)�-��Y�=W�+1��Y���v�#�_���ܠ|/�Oܹ
�b�*��v!��;�����T���N�d�
��$��e�ڔ��dDr�Z̓�H�DlO �=���B�c
K(���I�t��/z�n�����tl(�B[E�z�Vt���5���u6�x�蚷��
���)p~zf��`�'M6�f�p���cȣ1Fz�l�ݚ���W��3C�Ч�>�y�WQ��@�����cɦ���\z~���r���h��p���A����-g�$��sW�3����aA\��D�D�f���Φh9�a�P��%!��Eސ~��;�{=�jD�@}Fo@{�!E���[��,���v�\����� �R�r|�FA���57_-#��v��Ce"��kA��uQ(C� ֞�5�q�dW��+%	��w0�I��9���fr�����ކX���W!f6��ʸ���0\����;� �l���x�����'^�&.�=M�}ol������h��m�I{$oء7挫y��*�p����B���G����/��D��C�x2�j�7]��9�V����;��
���܈Er�������B� �yk�mB`�S��t��x�o������g@�Q�wrغ��$q!Ƌ��v��)�%*���*�ЯPK�0�  c
  PK  ў,J               213.vec҇oMa ���ܪ�j�Y�R*1����mR	��Jk���v�"���J��������͓�wNޜ��sCH�C�"���ӒV��ML��v��Ӂ�t�39t�kLB7���=�I/zӇ���L�v�1�!%�a'��$�Q���1�e�@!��d�$I(ҩLc:3��,f3�f��c>X�"���I&,��`%�XM1%��������l��n�Ml��-le���Nv�;�����c?��J���!=����cz<f�j=�INq�3���mj��\����9W���u��Mnq�:�p�{6�����y�Sb�����%�x��ڼ��4�4��|��|���7��g��#��3������f�PK���d  �  PK  ў,J               214.p��{<�m��m6���0�伊r.��hC	�蠻J���e����sw�v&�[� ��^E$S��9������^����y������]���}���~?q��= ���@@ �����4��KI#$R��ɢed�*X9����ZUu�u���iꨫ��746177�4�ڱ�t�&3s��E@$��A�ee�Z�Z��u��4�ȅ�� B1��hJ����!P�!�D�H&ܗ  
�A��`0�h�d�a��Z&$����3���'�cs�Iѵ닮�7-�RRƫ����o0��ܲ�j��n2���a������=q�� �|�B(����1�q���i��Y����������~Mm݃��O��x-�m�ݯz^���޼� �86�u������y�h���?��za$^
C,{���00)-8�DEx+h�^���$��mB꘹~Q��u��t���.��4���"�'�����-������|yH�O��Qw�V��݈Pv�_�"t�&���:��n���G&��\�]��YON�;���%w�������P����/�?�~�j/���LW�Q�w}��<�^�������M��C+�u�xXSzI>��b�������[9	i���l��@�)dd�	��k.+`���\�2н�c�U���l��{}��(���@j��n�v�Qvl|�[�EY����͹1'��4j��2fv���p�S�.�lB.�OX���T;�8ʭg��+���(�����I2�(�/���I&"f�s����T��q�����p��%8�'�S~"����hK���#����
�:AJ�.�-���x�Ȍ������NI����o�����!�1�j��~#��1��V�HL�F3�J�I�=��Q��	�
@˿:�Ӄx�r�lU+�sGTG��gzX7�C�.���6쌐���]�~�B/G\��ȓtm��&����g5�X>Wm\���diN�η�/�3،{�e��.�B��\���Σm��q5~�I[+�_CF/w��*�r8��6�R�l�]�h����.�%����L!��m��Q��.2��R.�X��h�	������F�-��Q\�g�m�GZE�^��G̖#��܄.5ڄ�3�2̰͡�~�o
1<����B>����Ӛ!�{�L�?���vym�\tS��N��g�ĘY���{��X��,��	��kAav��e�'��<?���4�{6��Zt�-"�3���<S�SĭO�v2�t}?��/�bs�NW܎�tb�4�JZ�ڣ&���$T<��V �F⺊��zO��(G8|,�;��c�{���k����6�T��z�]C'�ځ��V�Y^	��)��N�
�w�`��-n��TF��ܡ<��ɛ-8���Z������l��W�G�n7O%���ӓ�mH�g+159�8N�$����;� 6��s�`h_�}��9����R�ql���r%�Y��D�({�"��S��s�XԽ����J8?e|r_`��|kO81�,���&�5�5Z��@��b��]q���P�jcz��o	�'�k.���#{�O31'|�>�'�/����]}�~[r]V��v^��^�u�=3t��H8S,l���udoֵ�4.���]
i?U�y.�t!�:Q+oL��ǬeP����U�O�D:������(6�h���ف�~���n_r��%�����<�x��V��#lf�$W�d.)6ǡ�N�5�m<�qu��>7�jΐ�F�Ib�[c�R��j��Zi��b�WK�N�/���5�n���@xa�&�@�0��Ў�ѦV�7�%�3�<+�4I��"Tk��&J~|�վ�v�s���#&�1�7QvH�Z���gc���q̏$�#K��q�Un��MEK�9Գ�*>z���F�,^:�{��tl� �"18}1>���h7'�N�2�r`yU��cc�]�r��="�$Rm�[��VM%S�V:e�7PK��c�  �
  PK  ў,J               214.vec҇oNQ����S��բFl	j����Ml[bKlb������$��G}�x���77'77"+��S@�Z�?�M�Rd��֧�4��iBӔE��R�f4�e���i���V�ўt���BW�ѝrzГ^��O���ZA?�3��b0C�e�c8#�(F3��Y�t<��$&3��L�jb��`&�����j�t>X�"���,c9+X�*V����c=ؘ��&���z�6ݞ
b��d��ݺ���c?Ra�C�G9�qNp��)=��r��\���f.�e�p�k\����[f������=��<J)���k�>�/y�k3o�-�x�>�G>�g����7g�s)�#ŏ,�O�_ֿ���PKpUE�a  �  PK  ў,J               215.i��g8�]ԯ����5�����!:CD/!�'�0J�#zA�QF�O�w�{ѻ0}����[��眵��v�{����-�4a	����������9@ '#�����`

rJ*Fj�7��� �\�Pn.vNNqA>1~NN!9a1	I����������Կ�QPPPݠb��f�����6B@GN�
䂈� b:"��^����?�/#"�����)(o\O����@ b))	��h��8@BGJ�+�F�`d��a�
K�#�W�le29�v���dfaec�yKPHXD&+'���qﾦ��������������������@��/�"�DFEǼ�MJNIMK����9����]RZU]S[W������������otl|brjzfv������������c,�������\D �����Ew�ELB"��ED���	t$���d�jF`{>�0rF�ļ�V
~i�C&�Jf���E�O��;���/���_�Y�
Dt�< �d�*_Bӽ�7�K��z0=�ի�eW�-J~�n�S��:�!�נ� |�8qY�ǟ �i����=�c&ȿAҬO}�iD�f�rW���`a��M^NlC
�6����<	_���t`�3�&:�W�'�T�Z���d�fY=���H]�%�y+�$�2��4)��p_C�_�Vck��6+��ѽv��>�R9c�Mq�c��"ļ���M.Ǌ����|��̶��������է��n�}�1�Փ����7�;H��e-[z=���W��`�c�!�]��Ёq,�����Hu׊��EG��q�b�CH�yH��OE����0�� ��l]u����I�d�9��V�K�J��#�	�PC��?�򏠗�������{�ܼh����w�Y-X��lě��k;��t݂��)�	���4������4d�3Djz�1�H�d�#�*�-_�Z'��Ѐj�9��+�	�6�?'�(�j��o#^�t��=�0���8��f�K���ֻ�[���B"
<L�l7x�-6)ʫ���n��]i?�GTS�q���i���kqJ^F!ݧ�N���d�yA�{����#&��`](C�c�+K5KJ��g:�+T�hVy�����n�+J�馤�uO���as����@~]~5��&�Ky������W�6_`���%�g�?��@Wh8v�K ���EF���d+�9�%�|%s]�g|ɼz�ʢ�mU<�38>�������h0n�'>jDz@q�l�H�S�ݮw�����
)�#��AU=�9}�^��>�(9�1����pH�=������i���j�_v�l�٤}i]�=���]b�M�U�h���j���;��]�J���T�{~�j�]�o�2�[���1͸dPa=��t2�:��ь�/��Eg��o�=G�T?��\�H%_Z[(n�9�;XF�l�+�a�FP���V�wʻ`��5��|�&.��F�MO��~rnM�����(�H�_T�v��d�߁��$"�2as�Td�J�����`��Z3�aH:Y9�f��1�Hg�!n:Z	�u�r|�k�_VY�C׼��E ;#��VJ��1�]}g�dJ����J7��$Iet|��)�A�S	�P:^��r�Y)�>��@|t�JC��|=�5�U�!���X��gX
-�CNki��ܾU�%tC���}t|�W�Wq컰W�~�=!��~ C�q��`��}uD�h�{��CK��H����]�T�d;X�[�!½@yG���k�wq�6�yx|�`�ٕF�Y��% �j?n�LH��M�xK}��*,�m��Ȃ'��X^qR��I\��Q�yaT�$E��,,\���+E[���S{�6���	��l$����2�bZ'e�䘮�L=�����p��]���$ev!��zm��ϤQ����";�H��������!'�~� L��Ȝ�NЕ�� �G"�&����r܎%��}���i�V�h�6�V4����	?����A������̗�b{��F�9�{�B���-��:�ݨB&���.��E͝����0�I&��lH<^jݾQ������S��W��d]LVl�ri�K�.̀nJE�D�d�_
m�ˉD0+����t&�X�)�d���ӫ&�J��Jy�Z�v��G�����E����������;OX�)u���_H�N	��&I�Y��t�F�#.0��=�����腅0l��O��u�ɚ",�D�?{���T�̖��3��|�$ԫ�;��h�{?y�=��/�u~lE ����
W�t��T�Q��f�Yg��|�����!�ů���هg���#��ɚ�w��������2�L�&���x˦������Q=�Q����#�Y�znMT&x���-�/~�`���& <���j$�6~z3$��q��QV�,����������"N��۽�����eΏ�N�T�'��h[�;.l���Ո�6�k�w����
�ޢ_�����)t��y��lx��������g�I���Z	 {�C��˯���s"Ԋ�QG�P��U����	�?g��i>�x����_���ΛA�(����Op������{����m=�d����RP�&��1�X3�ϱ�\����C}0b�-��z�K;�?��21���E��_&��mY��sb혧�F���e�z��q3I��R@\M\A� %W�6.��0�R�.j�.-����N��F����I��)Io�w~�������e7��WD����n�t'
��~Q�b�_���ޭ����2��g�����ū�^���[��6���)��-g9�K��{���s	5��OhCrB�'��̂�R{��jW,{{��I�Q��e�'iH/
$�bK�t�Z,�H�e�~0(�gm��o�U��*�~p=��H�V|�,ʣkH6�Ir��e��xSTC��@����o���J�+��_�ca���E��L{��⠃��g!�z�$|���Z`��y�~��IuR4υ�|�T�1Z���OjINMs�;�
&�gX��(_���uZ�	a�R�u��X�r���Gfg�s�1@�w.Ko�d�3����q�9��ul�ču2�C$�x뇺�)������e�ޜ%��5���
y�֞�:��5Xh��I�׸���)�h
Z$r��9�������I�6�a7J��4=��B���v�kK������^��bd��D�y͒���9��	))�3�1�^I�v)bN�5d[�"��~cj$:����lx�u����w�������	NQb�U��)X����P��]���ކ�Iz�y����q�/�sc�z���?5�7�6_/i�xCs�������?Q��;|���2��ȶF�o�(�+I#�*�U���DX�#������f�$K�nɾ\�dY����)����ߝo���l�m��s���� �q�I��w�?|n6��67(�dg1%?8��w�E����T]Zn�bR��{�i��<���3��|�?�^�w��,�5�Ys�h��I�1�v$�,�):\�OJi"�����>�'��9��k"(Q�)scONj\qŪ/�p��?|c?��U
�yЛ��wz�t-�]�R>�E}�骚NP�1��w�\h�eb�1�;-��5R�s���?�Z�㰸ۙ�,��]so5����<R��N�(�jt��֨N�I���v�?��쨥��� n-������=�\-ZC�_���p��|w%��C���Q��3����z
�9u�y��5e����ʫ���'�sg��ʻi�M1�=2��&ǆ�n0��i�\̥x��(�Ed�X��(,���5Jۜ�H�|��[W��:��e夛��������d��m~�AS�r�s�D���Ãc�C	�!���O]�"$��b�u�Ex�R�?0��~�����o���{��d?/���TP�2s>�L���m�������_n�.�`��EjL��s���oH:�v!Gb%t��UGx_�^�|Ov"pi��2N�Im�?g6 �2GNa��x�^]WJ��
�%��*�*ѹ�|b��ND�y�:_��*~I���I�*�>�����(��Y�7��sIQ�E���� ���:�GnU��;9Q1�5�_S�1U�G���4�gŝ	�sI�:b˷e���>�׮��c�R�au��VY����w���?O��kWhk�gzE�y���ś"z��(p$��P�"�0V`����Ȉ�'�����v�q�9������)p�J�7���@�TO&� #�����u>;ȑ�Wt�_��	sI�~ �ei��1f͉�IZ���<%��ME8ۜ��6ts�2�x��7��(��?A��>Z{������G}�;�a��[ڪWt#y�"��ף
��t0��|���({�6��S*��dܽv6%Z����*M�{�n2_"u�&#�<�b�M�>��c�k��s�q3�d�<n�"�a�&����$!��|Q9��{N�,��cU�R�=�X���`/�z��u�yz�f����b�������ll`���t�}R�3֓����;wu�9GS�A�Ent=���ZYq+��3�$A��26�C�j�Q��0bf�nߐP`Q������+��4��#9[Oq^��X���p�G�o9��_�1Rf}�Z���/����	F�n���RZ����W��Be\��.���br�~�m�u�Kqǔ�����#��,���[���}#���i��?��Z}g����H�i�P����|Prl���Kh�V����κa#�@�׊҉��w�̂�ڏ�^��ʍ_�G+��G����J�+�֭�,������|eA��vڑP?�d���_B?��-�*�!c6*7��qX�^�nRE[���J�8MP\�C�`
^�Cju1�I^G����`H��>�
������1P��Ғ���%=�{�WN+����QL\аb7�M)�i� `�_��A�.��~�:��Jrg�ł�Br��.��%���T;U/�E��m�f0�h�a���K)���^���MG�d���~����,F�i�J����L4��:�oD��%0Xwmr]�����M��JF2�W�_�0_Q+�LC�u����
�>�P��<o�<+��N�ǅM)MA&5/=�&�y3j���3���e��O ,CR�.������ߪ��W%�f6.�I�ꆎV{�]X���$\�zZ%i��8�"��c��
�BIg�+��NH���p
u��jh�2��e)bd�T��T�|#���|c�0�|/�RD/Utm�:|�R4 �@-�|��VaY�9���,|���d�3e��*ܩC}ׇ=ٱ�-���ɯ��p�Af�بٸDU6%��W�ѱo�1E?�C�9�]p7S����f���H��@oN�b���3�NT>왃�ǒAq���_V��c�#ݳ�ώV%���f�i�&F�/p�cE���rhf�6�7�j0;n�!3�;K�g�<�6wIf>${���# t�o�3�%-���7^>�T m�%Pf��e�@�wE�1��g_����$j�O���
�gADBGC�QIt0Trh
c�UY?��-UN(�������^�>��/��%���I���+�?�,��Z[�F͒��i|��e�V��jL�¦c��E�C��
0�D�^�C�����}zq�O-�c��AM�<,ڥ�[�)���Ս͛�i��Xq4:�# F�O����vbpb��/g�;����̘���c��B$A�u�3OnK�����x�5�n_����]=ن!�#�.I}y��3��(��.+m|?r�'�p�H�@*=m��^���h.A�����֠����ܫ%��a����>�:��L�9�Xύ�P���؂\����ѕ�U��O\�H��Q�9p	��<�J�!�^)���'A�^�)w���Ɋ��f�$�l�Q"OKK�Z����e�s|m�}�`D rtS�D�M��e+|v®5�@q��nU��%d��E�l��?�ob��%�����Mn�)��h��?��fV�v��Mݚ�U�ԓ��
�{��ǣ�Jbs4g]bk�,Oa�h��АccJ�=m��x�t����1���Z��O� �H�wPRdb�&GBa�7�t�����/.�v!6wi�č+�	�9�6GD�`��=ț��u:�î;(�/m�5$����b��*5䰠�g���7��(x��`u�!��ƿ�P��gڟ�Bϩ������*�myE��O��9�u����O�����r��Y��pԓoىX�r�@�W+���Z�KIۖ�r����CNd�:x}ql{TA7<.Fk�;���j�/����d���u��wFE��, �Z��sҘ�[��W��������\��\���e��Z.�:�(�H�J���Vl7�G�q�W�簱�hrP�W;~˙��K��>�G/�s��3��tG} Dw�R��Ĩ�](����%�;s��]w�Y�N�7��"J���L)�Gl4�L�R��:s ��~���P�"��̥��C ��|L�R	&5p 	��Z+6o�����a�H����3퉳x��w�0��#�I�'�+O �ٲ��dJ�,�[N�i:K챜x6�:�]m�_�<YW�=�������g�s�M=I���pI��f4���mK����0�]��_-?�C;�?��.A����%�-���E�G-�2���p3��h�E�*�� �@��)Lz��{<3E�]k�G�J�!_���\s��H_�>�u�kj��Ʀ�sj�>�aQh�����F����sϽ+W�ǜ���v��QI)�R���؏�������PG��G*:B��E̽8�-'*�J-��R�U��&��� �X���y���T�]7e�{��y��ݎNU� na���:��_��WK]QT4�y���P�v,���v;ll6 �e��DS�/�wEG�I�����Ksd��'��⩃[�?�,&ӈ��D��#�3�y�(!��)B#U|�b�,���yu�=��sJ������H�l!bD�]pv�h��?LS�{ӊ����ϸ끟��c`�:�����-̛�ϱ"�*�I��%W
���$� ���qW�d���_�f���l����1�K�<)�2��"� ��<���n�J�x-�ى,�*x<��.{>Q�J�jU�7�V�1�et�y7��/��*�Wd��<T���K�篅��Ҟ@��K��rX���U���(>������N���I�t0���٤y��;?Q��쑈)�A�xjTgVS�K�v�Qg��HV�D���P!�����h6'�M$�S�r51���5�{�0C�?,ˑ_۹�ڸe�ߙ�cc��=r�B�v�>?�/ykk�>�Ѳ�0*�[��_�1<ڍ�%��x�Qr���e!6����";d���@�c2y済@J�KN��㤳>��r��ԩ*�����g�ne��fN+~T����NU���E�(���6��+wV���D����$�����Ϣ�'�"�E�ҏ`E���HL�F5�/��e���b�b�<���ε�R�q)Jl7���,�>�����mF ��+^��޿b�|n�Ҍl��Y�-~���f>��I�W�ٲ�&�
~B��铌SV.eHw�jrJ~`&�-�D�,,�L��wf:�=��р��pyW~Zu�;!u���t��!�Ą�$�3����4��C�����4gr3	���]�xӆ;N�'��y��'�����<4m��JX��A������� PK���<a  �  PK  ў,J               216.p��yT�����=bH�HLX�!�J�[dQ�#AFQ�
a�@@� ꈚ��e_��EA@�aE";�Ȫ�4���T���}���{�=�w����_2l����@2  �.@2X �"�p8�@��rhYY�OR&����DU=�*EW�H�k����T�}&{�vl$!�H�,� 'G0P#����X���(�Ƃ$O ��N(�� � 0
�#�(Y��m�����PD�%� X����sb�)�x�،;�����]s����!QJ�	;�5wRiZچF��ML�X������s9|���oG������)��g��CB�.�G�'�/&&%s.s�df];v�ǿ���_PXTRZV^QYU]����iSs˳��=?����������_X\Z��iE�������za�^2��Ʉm�B�jt�������"�2��#�w9�)z��B)i�4�7�~5������ٿ����
@�A��c3`����!�C�-�	��%�N�����R��
5�_?��v(ן��SR��~�I~�]5�E ��v�r��*�W��Ѐ��o�q��|��܌Y�O���O悗�+��*�0y7���pe���x��I�;(�RK���f��zK)�Ump�*k�7�g���%���z�|~�8�ݐ��g���N;Q?�?���;���.h|��j�P������dgCO������f�D��X�Y�MY��N_�(��8�	x'K�k�Fk<�9��4��!�?��N~�j�8w?���t�vy���=|q^=��a��+ǭnO�퉒�EA҈1�#6'�Jn�:�@�6\���乺�@���fY���a9�_}�d��ج�B�i=�s���*�z�����?�ٓD���������u��u���{��6lU/�x�(�$��Z9��,�Y�����o�V��m��%4���3��#�W�6�o���^r�Ƌ۲��a�{,�Z�SYU:)��=�9��x煀m��O��3;��};�ԑ�:zKWX\+�_WL/(��:�X�LZ��HYh��g�3K%�_�w���"�ۿ4��ִ����1ی.K|�����#�=���u�|U�e7z��}H����̅T�
�(�<��Z�;q2��[ R?���cXj��g����({�-��S�ݨf
��@?�1���g��ٛI�����x'�+(�W�}rV1��[1�H#���I��C� hW<o�(�)�����%�eT�ZT�R���klP����G_��AJ�[�H���v���bcd�f�1��2����D���,%�_�f�D��ާ�$�S�[ß��/�j`��O� 6�'��N�C&8Y�M ��n�kV>�to����P��S���P]����5�+QQ��7�nYZ�������hi3�3����BX�7�r-b,~��.�X�MLTi��S(Ќ6K13��K���gu.\��W���7����<[H�Gc_��~dc�X�]��ti�	�R`۵��񱫘��o�=>o/��w��W}�]�CRQ��{n�X&��J� 35� �,3QUԾ�]��K��E��ƨfJ�%h`9���7Y�mH��<_L���w�8�aU�����L&��y%'�4ǔw���0��7����L \��%ׇ�~��"��&v4^�V� �4��]r�V+x٭�X/�����wo�V��rؤ�Sz,����pV�1��뙠�����r�{�,˘�8��]�R����Mr����n�4 �m�ݷ�[#�����+u��b�8��>&�̾U	�s�8�H�U�(��O�81(oS(I�k�ܴ�|�Q;s��o-)��]�צ�S�3�Mp�Y�
�����r��D�Y�2rYq;~N���X���&{��	! �q��f�lِeC��s���c�>�`���S�EG�y�����`��b$�PK��Q�  m
  PK  ў,J               216.vec҇�q��������[֏�e�M?���g+[��&�l��&�l�)�u�x�z���^]�uY12G
���JU�Q�65���C]�Q�4L)�5vބ�4�9-hI+Z�<�h[�ў�ґNt�]�FwzГ^�β�}�G0�AfHV��:��`$���<g��c<��$ʩ�2��u
S��tf0�Y�fs��|��E,f	K�e�����W�jְ6�c��g�ߤ�S1��V��l��d��c�W�����9�Q�cz����9�Y�ٜ�\���2W��5���Л�ʳ��w��=�����P��>�Y*�����6��5ox�;��|��̗��k!ŷH�=K��������PK�IA�`  �  PK  ў,J               217.p��{<�}�����jNՌ�Z�):�
[���������C7I19�B�Q�""B����hN�L2��r�H�^��'��y=�����{����s}e/d}�"k� !  � {	��

�"�@"�T0�*��*������t4��W�#��]C��&m\�ƀB�іM�S��3�Q��H���
NUG�k�9d� �"��
u
��@Y�\�'��?�@ap�"RIY��l �P
��`���y �����
�Y�`5��5E�Yq�A8�g�ɉA*-Y����_I$�ZM3ڰ��d�������z��urv����u����o��а#G����-6�t����Դ�3.]���^��{��[%wK��WT�\[W��(x������)z����_2 z�vxl|br���/�3s\  ���%��`Pb���[�����v�#x�.5Zcv�Zq�`�0�������^�͡� �s`1�ٿ�����@Ay�(��O�'�$��B�r2��Q���w\���L1;VYPGr��}��w�f����i�2�s�1a�j��KQ���{%���|�p�,:O�؃�')tH�S�u	�M啓��Yh*a��?�0父GLnᢍ���޽>
:q!q4��]�6~	����E�q� Ke��GTb��̪�|rtT�YRv~��rS����xh3Õ`���`d*/�~�y��������`�@S�E�����Y�#�&\ԉ۶0��F�>�#���}k�u��/H�/��1l�Λkn�Z�,����p��Z+�͈��k��˶6�M��eItlP��AA#S7�jװ�X3%?j>m�-�v� ̃����`�;1Lha_~�dnp����]�"���Q���=���:;:�`�1�	����0ls�/#��,�1)4Rpk�|Тa+W	ȵ",ҕ2ñ�Zlx�f���S�w��X���~�sGx
���2k��ȐV��I�M�4�AZ�4��??����<�ZN��,�o��F��娭M;�'}��u��b�2uXWц� ���[�w{*�6�Sz����߰#�PȀ�7ˀ�i���;��b���ة�Q6�w.�4��%GD�k��M��(���cڭ>^�� �c��	��$�t�~:af����4t,o�d����3RtN����2���	�W2��kF�u�4/��4����"�ސPb�1�D묶S��.�z��]7�㊩�>�#�;q5���U����Op�@l��^����Ֆ_���{V�Zu�e@<Oܿ����d레�Q���ςٗ���=8�RE��?��ar��0�h��ty.P��h����CT[���S�j"����7�+�^�Noťi��}��[x�?�-cg���`���������|h#VxS��tq��ԉ[�<�Z����^M��R�>�Z����9�C0�8Hn)����[֣���a�������%W�	$w�,Xĉ��v�$q[7�`Ѫ���'�E��;-e/I%��=U���I��V��_+,�EXs({8Hu}))be �e�`k8]{B���$-1���>����#r�k��W�蓇>r8��\&=�����ܳ�3d�i��ђ^C�+�g����2���4��kLI�%w)�|�O�Fsl3^���7���Mo�^��T�m',N82]��/f�I�{r�78��T�w7u �
�;�P���Ɯ��^�����|9'���t*�Ҥm�d�Wa�c�ަ8��X�V��ɦz��w�@�Q\�S������1%�Cc��<� �U��ߢ�R}�Bw�� S-<�im�f��b���P�ྵg�w[�Qu�O�m��vw]���x�I����|��'�{���x�
b���ʖ��	Zۦ�c!��7�k��PF&�]�\���D��I@����ז>K�^�x���t;�4��,��p4�p^��T��	�Ɛ�<ٓ;��^���m�V�Ё�����8�.#���^�mg�
t59�ReW���h�ˋ�Y�Ⱥ�PK���  �
  PK  ў,J               217.vec���Oq����__d�q��l�d�M6e+[�W6�d�M�q�&��?��������t>�_>'"+F�)�@5��NjR˦�֡.��O҈ƩM�zoFsZВrZњ6)��ڎ�t�#��L�ҍ���'��M�fe�O�3��b0C�0��:���b4c�8�gt"����2����J1Sg1�9�e�Y�B��%,e�����U��S�ѵ�c����Ml��آ[��v*ؑ��Sw��f��e�9�A�Cz�#��9�INٜ�3����E.q��^嚻_�����csW+�W��>�!U<�qJ�D����e!�W��76o����G>�/|�[�o|/��)~f)~�o���PKJ'��Y  �  PK  ў,J               218.p��{<���sa.Fú�ܒqo�ĸԨ�ń�q۰�.�)��\�\ֺ�쉑ȭ8��̆M�T�dIaȭ̎}���{��<����y}_���|�����8i��  �?� ���0a!8C �HF%"�����(�)�W��b��+�h�b�8C�Cx"���nt�D0��'v.!�JFTT���U&���o�p�P � `4��;EA�B�?�g����0�@�
��0C!BBP� )�P���2���$�,L�"�p#��z��]�����^�R�+Y9���8M�aC���	s����IkG�34g��Ϸ����w�rȕЫa�q��'$&1��13+;'7�Ut��nI齲�����7465?��|�����|>4<�}1695�}3�v����e���ǵ���. �+�#Z��B!P��S��
)�%�Qag/J�n�1���������ϐ���jK;h��5�����O�s�(H0< ��8VZW �E"�~�� ��\鯅���~�!�&"�͌U�s���Y�sn��)-��ƹ�ܲ�0��:��/;���9�bj&!q�����
��ģ���(l��.��VU�'��W.RR��6Ʃ%R780\g��d*]���b�d���8�#�:| [�C������q���7�ɟR^
�Y/DX�z��#�_Z�P��G�W�d�_��VL"�8��2�q�Rr)9i�Q+�|��i>��w����M����hv�0�~YdiK�JǱ*��_�fIĽ��J��9���5��Y+ޛ�0��*ä��2Ed׍s�'�ny��5AUS0Np�	����D�{�wzu��da���6�r-��ήcs&*fLt��i�{��3�t/�]11��+�R�v\�Dzx*~�<����u�%����2s�j��Q���h����ٔ8�[�Ցѡ�4�j��!J�R0��]s���f��S6�##�DӸ|�["v8�F����6����)��+zӫ���Z֦X�W�$�,.r/C{ʺ���Ր"X�c��Ə[]ͭ2c���X�2�gFsL�9�M�lBMD����"X슢���W��4r黭�G.���w���U���mW�G��ؖ䐥ԑ�H;C�O�����<�5�y
�aWWVO��s���]�7F�EDY��g?��S&u]=���(�zkQt��I��i��"2�~�����T*�t�������W޸x���}�6P\�+?�� k�b���e���&��������n|�.��H���[�f��f�2���c;�8��I1w�~ef�6癞yk}WƸ�����9y�����$���/���9;�7��"5Xe�u��)�����	��[�𼕯/\*��7kmIYHJ�_������D��O�Z���
�4�<X�3$LW'hh�Xj���GNKS�#���G��Þ_U���řF���!<l�}傤B��91{��}k_3]R�n�.O!ú�O���bi\�l�A��"�V�g�.5ZI�R:�$�>�}H\���^e�yq`NT�q�	C�ٓˎe����>J�����n\11��#m&�.,�'�*��M���X��4��P{z�H�ɍ���A�5���(�s���0*�v��Hj�3�ԉ�>��/�;T:�|,=e��y��9��}T�.G|<J��V�{Z]ex\W�NZ��Ό����9���zв�y� �:ڌ��㝣;���%��Đ��5�����ټt{V�v�P�7~U99�����X_=��M�Ѩ����fa���,�-�:��b�CV�����E�5��`XH��pb1ޭC�����z�v&P�6��d8a�\i<�o7�L�2j��_�QW�3!uOI���r�ac�?�׺���)�[K�4�O����ё�`�#)NY>s8f#3={�Rqa�5�x��1�j,W�ܫ�sg{�U���9�k�$N�}�l�<v���C{y�B�ca� ��%Ǌ�_�PKM֏�  �
  PK  ў,J               218.vec���Oq�����{���le�&��-����l��&�l��&{��G����=?�������"�(���_�P�jT���5�Em�P�zԧA*FC�F΍iBS�ќ��Uʣ���-�hO:҉�t�+��Nzҋ�Y!�h_�џd�b3T�1��d�Cy��X�x&0�ILf
S�bL���`&����2��,`!�X������+c��b5kX�:ֳ!�c�nb3[�ʶT�u;+�إ���^��?��=�!s���8'lN�)Ns����<�hsI/s���U��unp�[���w���}�G<N)��S�����W��76o����G>�/|�,Ʒ,��ʊ�Q��g�����{�ǝ���?PK�q�m_  �  PK  ў,J               219.p��wT�Y��/=�0�&�PE@��b��Cɀ�����p��E���H�"�b4�R"�!@�2*�(A欻�̀�g�;���;��߹����+� YG�# B  /`�� �$�B"�h4JB
+-%))�	#/�U�������7kjo�0�TV�1�50"����i[ؘ���MH�I@4-%)���Ƒԕ�I�s��r(�(�� D�ʁ+<@M�N8�G ���HZBR|�B��P(��a0�n�x���1�D;��g R#KJ�.Diڗ6(кf��D$�%7�6��ut�LL���[X:�8:9S]���޵�g������!��FF;�r:5-��Y:���K��\��e�(�����w��W<��VU76�7����w�{z����GF��'&��_Ͻ��q�����@���^rb/�!W�@H��9\����y"��5HI(�}vaiZӘ6�p �KBQ�dx�ܪ�f�&����G�^�*���jVV2]� ��}�U#�k(�gWپ��J���O����*6�Q_��;k�����'3��ksO�k1#��Bi�z~]玖��L�~�Ě�cd�F�`�i;|�fk(<�N����!��s"����Ғ�����D�6ձ��3G� Nv��C�q��AAL1�����G�1���]uP 5�q��ȽM�R
�ÈE��h��Mڹ�[�FpU�«E�<E�zA䈫�p�񷱒�U!Zia	.þ�*�XJ
�u-3�u5Iz��	e�
�~��A5?�o�Ņ��{̜��h[���kw�E/�_�2:yF~7Yɾ��K.leD�k$
_���!�Z2s��4΂^�O	9E��C{��n�6�(�K���j�)���y&��qn��*���#'øq��G����g8+�*2�=�yJ6���xR�k��\���7��<T����&�#��FF!4?��D�>q)t/ETi�[[��Ke�}���[?o~2/��=s�L�8N�i�ƢМ�w�A�������ց���S^NA.���5�X/��'���Cmͽ�U�ĸ�;��R�r��Q�� �>+VA{�= X��K���x}L�b�]�~��%vn�s%����''�ߴqF���1����]�[�Ĕ�`r�#�o?6(�.�<g�g�暭��Wi&���T$I<Z�b�H.��̋E�T5��w�o_���� �x�uw�h��b^�F�Ȳ�,\:ҹ� ���t��.������g�[#",6M/�F�f?�{5��â�2��S�V����=��6�|�Fn���[��#v��zc�3�О��KH����/��I��e��T��r��b�z�f��X�.p��#��P�s������,Zq�JO lL9� ��j���A'�ꂸXX�'X�8i�o���-�>�ƺ�1���Ә�����L�2�����6�� �9�XpM%��?�kcp����J��3/�N�_e��&٢���3B�\�(:|�S[k���u�����QZ�vB@�7�^����X��jR.Q�5Z�kNp�R�*s��E�K[�+*�`�<�Y��_	������ˡ�	_���)�&��To���3ב�#�f`Y�W�R�Ls�6��g�o\���d���w�*UK�!�X���r�צ�N��̻Y�� (]�|�Ss�f��d�3���®?�$� ���s�%O�1�?4^��9�3��&fcv�~٢^2��.�5��9<Ţ�������[?/���Y��O�PxǇ�p�)+.U�@~�Sf؏��{��]u�wο";�GC�}')�X�⶗���K��9�
��>h�8�hR��V���b�ڤE.��_�L"�<�ʼ���PT5��F|����`O�8�?�5����f��4=gu�/>��G���A�]v*ǚWr{K��tsOf�ȗ��o��`�C���/��*�g�s?-�FHш�����4w&)e��F֨k�q3�r#0E���>KWQ���{R<Aq�ȕ�PKm�  �
  PK  ў,J               219.vec·�Nq���y���k�2.ʖM6�v6e+�l��&�l��&{��G���y���}ƧsNDV��@	U��*ըN��Z��ԡ.eԣ>Re4�k�1MhJ3�ӂ���5m|���ӎ�t�#��L�ҍ���gV�^ڛ>����@eY�!e��HF1ڦB�0�q�g���St*Ә�f2����9�e�Y�By�X���ey1��
V��լI�X��X��A7���lak*�m���y��]�f{�g�_p�C�G9�q�z�S��g9�y.�\�K\.�qE�r����f������]�q�<�QJ�X��g<�w��W��y�oy�{>�O|���b|�R|��%)~D����<~�'�PK��n*\  �  PK  ў,J               220.i��eT\��g���R��n�nB�	i�A����J�!�S��!��j(A�����]o|����Η��9���^��on��t4�5 @<  x7 �� 5 1��������Q����?����ca��023�q=�e��df����� ��*ʈ)<��� 			99�;3����n���@e@>��Għ���w�$�� �% >!�����Ρ� ���G�OHH@pg���	i�EU�h�^�8|�Ģҋ�9U�{�'�����IH�?`x������/ !)%-#+��D]CSK[�����������������@`Pp��И��q�	�32���������������������������c 184<5=3;7����{�������;�{�>;���\����[�G.�;.<|п\@���	�E�hT�@/|i9Ģ��TӋ�{H8ō���&I�sI��>��?������������ ������S ��&~y�=zB���?#���gZg%q�L�A�d��+����Y�3jR#L����	��w��C�B+��St%y�S���[���W��)o/m+us�g��Ko�~^ji)-2�N�WY��H椨B����$�~��� r��0����F���V��kI��!�b��.�'
�O�A���q��:�����&��G�J�,��P��ՆF���L�{�#̀�E��77�}��/,5e��x2;�^k���$҉����t�L\�0Vo���)Z�I­@O�,�[ݼ]�N�3�TQjP}H�v(k���ې�XVk�O�ۦ�k�R��-���,�zπ)�s MD�N��&l��i��r�,y+���QniAfHE@���G^� ��
7ʹ+����g�u�H�侫 Y���so��yB�n:k-��x��������zQ�G����Xf&�I^��J��pQ�><:\T�� 뗈��M$K�lr���$9fv��5
ڶ�o2�L�����y�������]���$ɩ��d�������s����6O��=ݕ%����]�j�	����*�xoe"'ǂ�-��:��`Jox*x�Y�7�Ķ*�'����?�؉	�\؂�b�:5M�Έ�ɚ�{�vI��*l�J[,ާ�#QX����9�m�q��o�oFR���1��F5�N�%�@�8G��d�qoX�[�|�6(�,3�Rn��g�-�*� /}���6=���9�γhO���g�&tޙ���t�;Y��
�{+��n�n>��m^a-gĐd�U&`��;!Ɏ�3�ň~��!١iU��g�?���������*�%�r��	h����B��F�P�/ئk�6���˹���-�!�	<Y�� 	�nCwV4��I��ɟ�(��u�J��z_b�ū��tS��z��V�8�idw�E@���W��88�� g H����mu֢ԩVF���
�K��r�v-�TY՟QPC��"�'�heT��o��_�˲�;�y�U�LT2����d�⃽����T:���ғ*����5.�=������OMPН~C�@I���D�kg��9���<d�8֬!��4��d�`��0ɴ�H������ƺ��=�%\���A\6��c��-��-$ ��P���`R��:?�u��cg$|ԏ��Q�g��Ԏ�|���ِx�e�����Z܃L�2ǅ��Y��r��Z��~��5�t_m�0��$&�W&R����z0�*��^B�D��Bzu�p����;�ʿD1댠=�OyR�Ѽ��}�)b����}�>]�q�}�A����>7�v2O�j�M�3|��|*��E':d9���G�� O�y�.Ơ���z.Ϩe&o'���rgtt��~��ah=���F�����>vX�f�R�nZg<L�&��k�5�M�&���n�!�"Q��i�yd��Y/�`��nJ'B,�ıUY!�iO*��N
�c&ZԷ�w��a�ώ���B�lc�i�'�7{t'��g��_�U�����O���r��E�_>0~;�����X�K����b�͡��уJ.���ƣy��>�88Y�fT�h���!�ʂʞt�٨1�G$���+�%X��� ��ō5��j�����,������'IU�K�+�7ӭ3���=��z��[4���e�+����4�j�}���M961���s{(��;��'����K�����Id8���-��QY��]��'~Զ@�`:��;rk��J,�I��=}{a���P��vT�M��e������NiR�~�iE�E�����obo�[�{?�9d����s!����Щ����GE�w^���C>��o"UnMQ�j�bb̆%>��\q�X15�����Mv_��fW�7��D
+�8nu<�V��Mt���Y���`��?��	=��������3���aw6c;�߮(��-��3�f~^B=��g����x��+��Շ%)�a�R����X5�_φ��\�u�:��ȉ��w �Vך�\`2�eZ��h��V`C
��-U�x~H���z���)��xpjHGP��N5��R��q�v��Ȁ�� ����f;un��أ��]������T�U�[@*���tُ&	D4p9���{O�Rt!�����y�� �܂�Ϫ�+�B[�f��G��)>�1G��~�%�u��O?[��G/%!w����q�BS3�R��*[iJ'x�t��1��㋞�t�3�%���d����7��8%�*j�~{c�0�z�K����zb�������U-$ʪ��*C���C0P�Zh�/`�aҳɭ�ى����xJg۬ަp��KG��P��������:��N��������^�&D>ܣc١�mv���w�:��p�p��
xʴoĒh��aK;���XQ	�Ȟ�j�T�S)n|�wVJ1��dB?���9WV���	$�%��-E��u.Y�S/�ɶ�6���
�[�0�<����7I���;[5w�ε0~X[�I�ǟ�Ms�3ű�n�8�1:ǿ�sv�g�/d ��d`nrA�]KW���q��ž��h��J�AMA9f���Q� ��P�z����u���n�*��>j�JzU6�|�FJ7D[�B}�k م���a� ��pis������<���?q���eۯi�~ӬU�e�����G���"���q��IEͦ�ӊTS���k^�n'�ʑTS��>R�F�E�V��������ݸ~ϧ~m��Z�T%�F��z��(����?g��`�z��n���\�尦ˆ�"+�Z�"2�E�iR�d�,��]��~����3+r�l���[�]���뗍��2�'=��&�q?�-Ix9�H&�w>�heΆ�MN��Qn�*0)+��bf���L�<��B�h1P9����n3ܞN�t=Y�*��u�)�#?�\��:�4�#s��(���&1�MU�7�¦0�̙?8��6�_s�W��9��=���e_x��T΄ic�Xh*�as;ߵhU3=�F��6��7���8�1�9�1w1���p��6蒀e�]��E�v88�Ey�o@f��,羑�h+Y���n�*_�h�Զ��1��ei���6YY���YPV���&jXH��L/W��R��g�<qek�����Μ'ޅ����L���M�;����1��Y�~����t�2��䳡	?�Z���W5+G_��<x9�5� ��5���
�6lͼ��5�+sz�}#ſĉ�6�A���[ J�L&�����M�����	pnq"�V���>���VW�i�S�+I+�J�	\����튣�Bγ6��"���f�󟾤����f�A��o&\#)wJ��=+�F5v?κ��Ur8�7)ײ5L�*a�iB'5dF���h��Jy�-ظ��(�ԇ�t�bC�tX�"M�bT�HW�G�\��&��V�h���y��sqJ�Qd�'�<$�1������� xAoWkU�q�$>��(q���\!�� C��()�@0��^���R��&��/�	�o��T=ՒΆcl�ɰ̜�]Ȯ�N#E&����k���\���c0�>@��"�E{I.���zc[���?�U#��k)(�-���IF��:~���������3y�%@�ٖ=���Z.,�k�:'��E���rƿ2wu������}Dr1T}E���4	�z��):�EGVx�Y����XΓ"����|Àqԯ�f���H�����.��']�2S#D/g]~Z�2�\[��Ld��c�<O��f��𵰭Z>¨����^A�T�VZ�v�(j�3S����_�;�8���O�k�Oq��e�mj,Ы�����W��Xe��5E�!�Oe�x�R�ͻ��7�im�³��%-��`H�wx��$Ƕ��79�Q+s&)�Bӿ}���2��~�.�Py���0Ku5�J��9d���a���?͹��䉆��7m�4��P!򕫿n&�)�;q�7��n
u(��c"�"7�6��5�,��Qn ���]��1�R���:�4ձ�i��Bzi�>�s{�!lԺ��n(v6fڥ�=�m���R�.Wp��T��T��r_c����?缠h2ZDTY�;lB�ی�k�~"�mc��ʚmy�]�5�r\��#���[�{�ǤZ{�ˑ0�U9D�	#F����h6�O�S!&��#@]��{r��NA�K!���UͳF��)څ�O
f�6u�wE��ŝL��:�Sn�Cf[�_Ġ����()<.��KM���~����]]���y��;�!�7c��Q���jf�P�ݯ�(ބW�R��u�._P�G�7'�6:S�o���e 11��yX�ϱ��׭RW��|�b�4T�
�ds�]�a��>�I�$���6iW�N�̂ `j_�Y���<��e��fΘ���l�DU�@ù�ᗂJd��d��/���<����:5*F|����(�rJ���/c1ـ��ݧ��!i�[vTn�J�!@�($&C�������my|�g#�J�v�2k:��T��vl�� v����=N?~�	���-���k��+9Yas����b���W�WCR���ā&�g���|��=���z|�3�^��8JV�e�q�~��A��4�R%RhԖ����;�bL�_[͑�n&&���Y{+X������:O���4���/���^H-EC��"n��<�P�uW��O��X\����O�.oե�x3B]��bY�����TQ�
�8w��<�!��4�fzB�O�|&񿬽dX���l�o�k�m��z�&/m	/�
�;/^����ٛ<�~+]���;�����7sPe�֗�2I�I�D}j�DbD���k��9S|13es�C�΃솴I<�uT+��c�zP�!)l�";lIs ��}�_�ǭlr�Ų����i��ٯh�%��cj��Ά$���9'ζ2�i��H~�<��!/kTk��_��������v��J����}@jЬG�\�݊}��)���r����N�.Մ���|�C?��f�4?m��.����]E���tU#u:�q�L��+C�y!���4�AJ�T(��R����jE�8k:��ܵ�~�����������RGߞ�����K�ӭ��>���$,��R�r�m��1\���wؾ(� 3�F��:��La��.g����ue��7��t@c���#6��#j=w�.X�"�Ww������'�Pnf��'<?�D?nzW˸L5�z�;��>�}X�=D���^��ӳ�궿��u�hO�XP��3_��*�}�o{���V���6�ފ�h�<B}AO��x\!���G�@uy�o���IOXe�Lo�<���k�_9[{�'�E),�/p?Z*zi��[|��������sQ���C�v/���)�[D��_]R
���Ί�?�\θ��\M/B}�ڹ��O*�zFMV�r3�-$���P�e&�t��&9�2����н�yO(Ȭ~T2�l���ľGDDu������uR
 ь�sEk�>�j��p`����3B� +���1k�����<	�"@�d(����Bq�*[�M1��f�1e��_WPk��t-��E�}��鸓�IAN�m�o&���̗�q.S�Q��{ݠ���s����t�՜E��@1��)kdJL����6-E���w[R+1bP]9�<~���I��L=��f�]~�X�;ܝW��*/=��'#�?�d�[֒_��9��7"PP�s�52�@;�P���������!%\e������+[��t�E=7�������Du/�5%�7�r�*�O�� ���$�
�rj����u���Lݷ��~U~i�{D��B��0S�o����b�/J��MS]Rb,�ʸ�2�[j�G��w�_��I\r�:$�=��C�,��x<~Z�OiΨ�3L��e��Q��b5ʐ:͹�^�����S�,�Ix;xX�vR�]yk�Nk�$���	ɢ��%����tFw�j���$2��A�墴A�]�G�Ldk��hL�\r�\��{�my�_'��b�Z����X�(˶?Q��H�ϱ����R��x�����I�g��
��F��ʜA�������C��+��6���@$�[Ư���Jc,���+�%V��!b/��|X@���̣m#�����H�<>��O�\؁�F�\����V{K����I�����7P�.<�q$�e/���ȧP���M[�>O�v�%�~RM�+�+����:36-�6Q�[i͍���YK��f��{5�U�DxQ�Fv�	aF�(��Ǝ�Ģu���������cx��]����h�c��	�S �1�>�V����v�^��ߵ"�z� q1E� ��@��o+��L{kt�I���]��k��>���Ɔ�b������$t�_����q/��;�����쑿�����Z�#�K���,/��'��p}�{6_���QE��X����_���O�G�U��)�]�Lh��H���S���/P�nm?�e�.�ZbL��9qȢUN]����p�'�̳��Ü�!�������d����7�����`ŧ�����T�>PV93nK�y�2�F����""��~�k?�1闧l ک<Z�K(�_�ūon�K��Um�=P�-���~a!K����r�au��pP�g��c�Ugʏ�#�i�8�&ۨ�TrE�C/,;��?�|��f���2'3|�f��LG<tS�f*��+=�y���M�ð�d=�*���sgL(}=���G�{�"q�>X�U�&";Vd_�<.Q��L�a��ͽܿ���O�{V\��l��m����W.I2�]Y��F����:�%�� �e��Wt´��QI�D��d�Q	��r%C����VVT���:>��8��l���A1��dZQD\�`���&�"�p�gE��/5�bъ(q��)P�{�/�E)�4EE��Xϟ_���/��\e&<�|��?*=i�ȹ";'c�TZ��Ŝ:h;�3�82 �\p�.O����ɓU �E�@�鉃]Y'q����+��l璝n<u�L�x�g��q�԰S��W��5g�l��$��ǔw ։�[+Z���w�q�B�C\S��n���!�����i$�2�Y���L g˖
n2u�p_�����S֜��#������]`�h�r"W�O��Wh�u�Z� 8��_�����+dd�>{׽+>��8o��wc=�Y�G����� h��򢒒���� PK�j��D  �  PK  ў,J               221.p��gT�Y��)��	BM��$��L!������0�"�QZh�HU�"m'�T�&%���&�4iJS�B6x��/+������ӽ�9�����+�[-�� 0 �D>Ȁ��8L\L����҈-�RRҊ��d�h�eeU��U��4��1?���c��F<n����u���Fnقĩ)����6 r pR�r �H��E}������!P1q�\RJ��j+ A `(DL
͆�������D|���@�"�r%4L���i�z����Rq�N-m���ួ?����(�,Z>b���t��݃��u�ۇ|&�,+*:&6�B<'9%5-���ky����w���������ڦ��m�|���޾�g#�c��_O����_X\z�aye��:���տ�q��P���Y_ SÊ˛Pan�m�H	�iRnY#\��nN���O$�k��_G�J�����'�?���5 HC@�Ã�D`��!��v7�6�W�N�2gki�b˄A~R�>��cKBg1��G]?��@thдg�����F.N�Ua^}���~����㦋��J�����i�:l�����J֨ANh�;��������MÞ:4����f������K���!�̢��EUS������`z��\�Ǩa�@P)����j��H��3� 5��7���
�ޝ�bHg��7�8n�\1��}T�E4�ꭈm6β�$ۻ%���96�.f8�^�t��#p��<��#Q0l��k���� 
bT��w�j���vю�����59�������ce{�4���=��{}����ޯ�%6Ty,Q)N�s��9.^e�Tۀn�	��M���ӂ�"g��rˎ��d%�?1��v����x+*��h�J</�S�Q�_��&�t��I��5ĩ�g��t%���x����׮g��Kh��Üמ�'�m�7q0�0�<��&ϓ�J�\�Bߣ��医V=}�a�F��)Q�>��$;�mDrЦ�u���A=T��� �|�5�֝=b�k����KaWK��ϗ4����JL/��U��Ǻ.r�GSMH�8�k��(�5#)�k��刦϶��+gV�e[�a��7W��/�3*f'�jZ!��Ⴚ37�{�?_z�F����,��!�r��$��|��B��l����=-���s����C����K��[��q��C�	�jW���������^Ͻ~vJ�E�XX1��:�`���4�RlE�~��dn9`jU�r;�rN�lXc�B�),mз�=�2X�y��r�bL@�N?���|��m{3Ӊ��\�"��ؾ���k߈�ws!YZ��3��_ʭbA,�r�M�j��mc�c�:������7˟J�Z����@h����qt���\75�W� �,�R�W��^o��b�elÇ7��dd�$5L��Z�����%r0Ez���!Yz޻q�i����8I�54la~I�����,$g���GE�d���Zf�����M��&�e��:xun�XA�/�*�ZJH��5��}_K`�>�oU�#4�5����B ���7[_W�7:����q΃ǯ�Ss+���S�!��=Wr�v�3��*�/�;o��M�=y��D0s����R�1���Z9���I���]��#��C^c��$��%��C���KSA��!���⢻���`1n��F/��B �w�Qj/�%�"��n�0C���
�Hn���:B�ݖ,��Ay~~�j}W�1�qָ9��uU�tY8co4��X��Q燲L���}��±�n=N�Qk�	�>��og��>�U��E����fhio�N�e��Ѕoh�����o��)�C��	�P<�� �-ۭ܇
�Q���-NϭX�?Y��� 
*J�Bz�������L�{��	��PK�r3��  @
  PK  ў,J               221.vecχ��a���}����V�l��&���M6�d�M6�d������yo���>wwߞ�'"�E�PJ��T���bSU�Q�Ԥ��C��7���wn@Cј&4��iAKZњ6����@G:љ.t��S�ړ^��}�G��AfC�p:BG��Q:�1�e��D&��S��4�3���b6s��<泀�,b1KXZ(�2]�
V��U�:�X�kYg�^7��MlfK.������B�Н�b7{�k�O�s���0G8�1��z����4g8�9��\Ћ\J���W��5�s#縩���J����y�C�G��'<�Ͻ���k}�[��|�����%��Z,�7��9~D���~��\�?9�PK��� ^  �  PK  ў,J               222.p��y<���cv&5̈�2��\�,�3c;9����:!�I�E8�]Ӑ%۹����c�ص(c;���2Ha�0�e�;��n�8����y��z���y�������A1��h�`��  $��P �Ap8�DH�0[P22(%9�����
NY�������TV&�����[���'��D"Q2(�-[�ԕՍ��7h���4 )4��9���P���@R`G �e$j�R 0X
�B!��%�< AC���`�4/�F0�(:� �i]����A����Vخ��۩�C��e�����|/ņjkg��x��+��;w��'��O�=w�B�Ű�ظ��Ĥ+���Y�9�?��n޺]\Rz��ں���G-�ֶ����{���s_�=�����������ϋK��^  �G�G/��K
C��^ ���hT�&gE�{�kE#0�iU��$�X�i-�ѝs�j��9�����b��z	�� Ix`4@>4ؗ�7A���7T�����S*��]���~�`�!:����
դ3}߀�[,�E.��	&�`3	����9�Ui�'3�� �a?���B��J&���q�Q�^���bY���maF�D%펿��#o`gP��E��c�wI,и�<��/z�h��N�R��i���'a�焥�y��l&�%f�R���m7P��O��~6�I
��4̩��q9��Nq1t�Dε�"A�#�];@�iҕ#Z��:*X�fp6c-���V�d�p�������gE%��F$�Z��YB��J{қ�lV��Q|F�x�h��~���v~��t6�����^+�D�8,2.iF&$���E�I���Nm�+wT�!̍�ó�d���{ϯc�\bT�ٲ?��?�1�1��i�\%|j���f3w�ahT`#B�2q񸅠�6��ϲ�-��N|4+�+G�LF^���cJ¬�,���}^��笤���j�fE�m �:F�#b�MR(8}�,"f7dD\��&�V�<�>�W�, _M�WV��Γ�i�Iӏ]hT�G�\Ɩ,��$�D��:�W���˸	�{ܴ��<�UM�����8Cv����@���@�t��oYQ��r��Ƚf��-b��G��Ԍw}�����\�r1`�b'��NӲ���ռ k���*��A*n��H�|�	�n"�}��2�GH�z ���QI�ܤ3
+���;uoWj͹�k���Q����$���TXw�Ӱ�ĵ=��aۦ�:krY,E ���ř_h/`�#���L��~{�}�p
&�d�Sra���V9enhE+��Mh�̧Ճ3!���)�1�L�+�L;w��+���:^G��5��sGC��;��jS���ɗ�&���������Aұ˳SGC�uߵ�[?����$�Z�<��o��V��~�&m)%2�m6�&Z���$P`F�BE5k]�nRr��1b��v���9�)矊:b>Ӱ����6 44�x�1�F�����
��谴J���/Vh���;ۿ���P��+l�\��sq�;����h��j�wV�y�P��N^T&�צ��'ɳ�}�4L��iB��v�0����k-��l�狔���M�0��c�U���7����N3���Ɵ&-)���}�O�����W^�y0�'�͝�5.��l��l�ݓ�@_Y�ñ4��ж]�� ���k�lS��r%/N�W�tVv�˃�NE����k����Q���g�Px�l��udX���fnl��4F�Ko����fN9���)�b���QN)�?p�������o8��$��G���6��P1Λu),��:�y,26m�t���S}�3�Հ� |���v}%զ]7b=
ΫQ1.���ſ#(��Nx����)����N#��Sʥ}�y;���ny�v��ڥC���Z��D� �J�Xk����PK�խ�}  2
  PK  ў,J               222.vec����Q����{]d�]��e�M��M��&�l��&�l��^����������tz�t"��Ȝ%T��Ke�P�j6յ5�Em�P�z�O�����{#ӄ�4�9-hI+Zӆ���=�H':Ӆ�t�;=�e�K{Ӈ���?� ��:��c8#�(F۔��2��L`"���U���4�3���b6s��<泀�,b1KXʲ<�庂����uM*�Z]�z���Mlf[Sil���(�Sw��=�e��~=�Aq�#��mN�INq�3���`sQ/q9��^�׹�͔���N^��z��<�!�l���缈<^�+^ۼѷ��=��'>�X_�ߊ��^,�%)~F�_�~����PKY�>�\  �  PK  ў,J               223.p��{<�k�s�aø�6�Lt13�dH��ʰ��U��%�2$�a\&d"�\�mʭi�B#��㒐ck�Q'�QZ�3z��gcw_�}^�����|�����>�a�K@i���#  H� �(�  �p�D (R�S@�ˣ5�U08-=]-mm��[	�������6�������;���o���W/�P(�<ZCAA���Ɠ�됶X$�(�� 0������N�k ���H����@� A `(�Be��d� SƓ��*�c��8r"�i������)��l��������1������;K+���h���8�u��!w��G����O����bEǜ�MJ椤��s/��^λr�Z>�����Jp��������{G���E]O���~y>����^�O�y;;7� Y��i��*�����+�C�(b��^=����$��=q촊9���+��2��~P�&���|�hv�+������ ��s �����"���:"X�����\��l�g9\�������_���29���6������6Y&~�����@.�Z�N������6�sهks�v��a����^ǷNCæ���EO�����ڎN��WՏ|�4rt ԐF�i�q{!��V��l�Tc�$&��s�B�S�0k�:�����w�����4�!4�����Vǻ����p��3�=̄�W��I��n�[�������^���W9Kh��đ�@�}�ΥΔ���0o��-Q��!��O-2���{�;�!���|.�� M�������7T���ȵ#���.�3qda�J�dwz��S�n�fcH�AV[3s�N���vkI�
׼�&
�ՠ��p���;9��$5������+ߨ'䒟�C�V����d��3���z��Q��fP�t�j$����=�<��Z�n�59��/���*��O��H�o���q�|ew�8�խ�μ�uSx�f�qS���:7ǌ�u�����F3s/ZI��!Me��c�W(����{@�C�������L?6��Tܰl���m��9{*X���6��:���^�в՛���خB�de�V��h��:!����Vm�:��'L��������_�t@r���� :�m�!���<� �߻���/�:j�F��#`QK��QR%����=ћS�z?��s�7�&ܵ�X���[h.��ӢGф��L�k�B�Wb����E���ы}��J�.��Pt��X<�e&<��o�ddZ�gخ�<­$��RyhX�ñ=8:���㰚q7K)�oRJ"�C$U�Z���q��{�=/.�@Y�z���3L���PH_�*��%��א�<�9 6{�R;��{`v�8�Y�*��4�ϙ�����4W����'��u���k�^b'1
ȳ�ѝo�1a_��'��ڮ����9�v���+Eb����q��=P���m��b��!���j������+�w���e?���G�Z����-3����m�C����A�-��%���`�_������j��q���,�nń�}��`�݊2���ˍ��������,e�z)���m��'���9+/�f��'.����cԃ�+�1�t;¼+U���	�ʷDGo>���Dͦ�F���N���H|]K��s�h�mG��M#{=�j�����"�^Tҝ�(���3<�g�L.��t��>��6l�^���´���Q�����u��ƿcR 
u|���7hL�-��ݔ��W���۔�ȫ�+�Bҧt���r�>���^z����=g����Ļ�i>��rO���X&�v����9�.��|),��!�m]jHo�~$�H��C�.���4�|��ӡ��9��l��a�juߩ=H����]�2k�46�'+���9NƧ
���M��)�%OPǨ����$�����J�#�PK�|i�  W
  PK  ў,J               223.vec��oNa���y��أv�H�"6�	j%��vb���&6��Mlbֈ�G���%'W>'�yNDV�'G���R��SǦ�֣>hH#ӄ��o��5�ޜ���iC)miG{��@G:љ.t��)�=�E�,}�/��� 2��ɲ���F2�ьa��8O��$&3��Lc:3��,f�[s����c>X�"�u	KY���r]�JV��5)ku�m6�F6��-lME�M�����b7{��>��z���0G8�1�ۜГ��4g8�9�s��^�;\ѫ\�:7��R�����gqW�q�<��c}�S��������6o�-�x�>R�'>�TǗ,�ך�
S|/H�#R��U�/�͟��PKI�K�_  �  PK  ў,J               224.p��y8����/H��� 3�2c-5�뉱/s�������'�D����r����H�,Q�҉Ld�D�"��#s�y������~~�����<�����~��.q?�ށi�@`  I>@�XH8�!
�DKce������e�*Ս*ee���QM���L1��٢ohh��e����\�fh���B����ddH�$��]�G 	� �@@j �`@�@UrN��U 0
�#�(��dC�z �@�P�JVc%� �#�[��Y�j�X�i�H�U�c�k�'u'�$
�ߠ�H��Ԣho242615�jm�`���;��{xzy�����}��q��GDFE�ğJH<�t���q�13+;GP�S��k�oܼ[v����AEe]}ÓƦ�ϚE��;^wvu��}�a�����ܯ��_Vt� �����0]`(E���#W6`�0�>\Β��*�fp��J�/}�"�\?�8amh���;��+��P�ׄ�����[�t� ���<��*)�8�h�G�Un�h5r��s��l�CT��&��ֵ� ]s}r��ig�����W��t
�b ����+/���1�XH�yjY�a�h�mc��y"s�O'�9��0�N(��VJm������\n
Ȳ�)����ۨ�f����x���F�D���5��]nVu�*n���p�:�M�p�Ay_�Qn*�X����һ:Bէ�&9�G�Iן�5�z �PM���Qa<˚��S�w��7Φ�^�)�5��T�E[�"���'�Ä�����Zt׃����w٣,E�.�dJ��%E�kO�(�7��}�y#
����;�v��[�7[,�\�5W<�`�)���P �Ňa;�Y���p�.��ZSI��1��k?�p��ڳ�G�},��w�Ϩ;��u-K�� 5��Ꮙb�w05l�K�z@CҺq-×��v=�]G���~]��n+��*¸�K���=�s�}R�Km���/|����?x�:�
x֝}���4������p�T>���{:�7��+R嗁{!
-� ���1G��db��[��g\��t��ܪ�P������1{M��[�4v�b���h��PX����i,�bՠ�
{��$^!��դ6�F��tc�fy�gѷ�So�
|�h��~7n���V4��Yy�'p��G���������Vn	Hhf:��x��oO~s�aN���M۫��l��9�`�rF�w�b��+�����56g�P˗?&ףr+vM.�U�zV�%�ӄ�c��y�F)�V�ȗo��҇G+Z�e'��#�/�	#Yc]9-؆�E/����l�%�������<� kM{���^2��=�h��-t�@�pjg�5��pl(�HE��W������=�1�����j_X+O�9���,	��̎�t�e�̼������\O�xe�R��qrZ/¹N��Im��a#(�j[rd`�tֺS�{�
�=������Y�h�b�Wc3�a?�\�㾨`/��NB������!�a��E�3s�'4�v`���h�m� []�q�	�YoL����@�����>���.ik:���e�qF:�������i+Z��a-y��ߘ�y&���t@�y�˔z��Ȧ>�k�b�X2�.�U��$�ﱹ���n膤V���L	�<c���qW�-����=�K�
��և���P�o}�X�;�� �{ӶRŀ� ;X��Nо����m�eY�����T��5�y�ǵ�7��/�_o�4��Dj��-�e����{�m��V��k���,x��r/���G���\.��Wh4y���|^sYx+�-�5����"b(�)=H��=�s��G�v)�y�;�=!q���\ɤ�0��e٭������OoG��ߌ��� Ǹ�,��������;q���P��56ft�}�:�후Vc�����R�'H7�l�N4�������J�u�/�:�?"��C��t��8�7���P�N����z��ݿPK_��`�  n
  PK  ў,J               224.vec��ˎQ���u{nd�]��e�M�le+�l��&�l��&{e�Q��>^�z�>�>�_�����@%��S�*T��Mu�AMjQ�:ԥ���h`�й�iBS�ќ���iC[�ўt���BW�ѝ��
�K{Ӈ���?Ƞ,��:��c8#�(Fg�:���c<��$&3��Lc:3��,f3��y�t>X�"���y�t9+X�*V�B�ѵ��Y���&6�%c�nc;;��.v���6�t?8�!s���9�'8�)Ns����9=osA/r���e��U�q��7���w�.����0�x��y�S��<��B_��浾�-�x�>�ϥ�����ZJ��{Y)~D����������?PK�l��^  �  PK  ў,J               225.i��g4�����,!k�������ނU�F�-ѣEXA"a� D�Qb��{��DY%:��{��^���]�����Ù3����33�	�<@���� ������LFJ�)(�)�詩nܠb���г1��٘YY9��x9n��be��+,"..畑���7	�*55L���S��m�V JN�d��n�P"���������?�/#"�����)(o�����@ b))	�_��_?@%��Q"�ӷ�����&�R���`0��-f���d�cb�����/ .!)%-#��@UM]CS�������������3'g���>��^��{�!<">!1)9�SjZNn^>����������KCc�϶��NlWw����n|brj�������������������ſ\D ����������D������� (	)���>�Ɠ�h9�r\v�
.1�=[�%#�����C���?"�?`��k
���޶���n��J!.��`�H������3N	Q%���g{}h\���59p}��ڪ˶���,	��p�֏ �>�\��9���cx�O��'�H$��Q	4��{::�X��Ә�s-)�-$e��3.�6W;@��vLz�t\+����Hͬ�t$�ڗ.5~�$�s�m�-�7U`RUdZ?V�Y�ͬKK��E�{�UH��W."#���_�Z��k�m.�r�9�&�dY�-Dڇ���W����ED�_���.mo_�}:���BA��!�Ɵ�i�}6r�J\����-�I�"&��%D�o������ nw��p��"g��H�V��F������!^"�����b�E����׵��-j�<�m�7H�k+Dx��o��{s�{6&e���>��x���� �@�]��߶x����	��(k@w�q��2is�&m<0���˴'��O4�Ψ�|5C�Z+!b�1��EV��t�����ǜ�y��2�X�x/�:��{��ҁ�ɧ��T���b����%�ֺ
m"��g1�&��ڟ�ܝ?=g^�NW�{1|+u5������em����dù=�-n`�q���u�[&�7��&ݱ�_o��Sأ{b��#���rhLy���2cU�����H ��P�ً#Ax%���3�[of5'v� ,��YȮ�a�Q��}�[��)L��wȹ��>�n���}X�-zBqaOB�y�l��H��!%w��5`�����H ��Z��ԟ�$6c���?���)Ç�'�_�}NՊ�x��ki3�c	/-�P"���#�A �C����L����D��t�E����n*E1+N�m�1��;4����E�o�\�8g6�1�]���._0��ܨ�H<�$�C�7�/�V��!F>�q�M�� �5+�;���e@��cGq
{h��ܧ��K���ܡ�#wus;ئ�����D��;TMu�!��T�_�7nV��w��E�M�.�DJWi7C�7"��<]X�bd�Fy�a�OsV��^*�"o�w�n)�ù�~2\8��HZ�K�x�*R�řW��MK݌W〟Z�u'�VcZ��r�qwy��d^�q�_$����ا6��ְ%<q��Lxt_o�o��-$B6��\����"��"z��F\,߁%�b��n�&K>�+O�<����v��dI�4(Y�>��@y��ͽ_��͜��;��n�]r ��FWA�H'��
��H��F���W߮"����B3���cn3v��D:�,�� �2C��_��{Ť����N>��2ȝ�F��K����,B��9���ft���,�j�=cu�����}�r��69�}��Ö<W�w��s�!�?����	IW�꺈�z�\�@6�<2\�f�E�CLT�x!_�L�! L����6O��]Z���������,Ud�[.�U/��k���7�?��i�ȸ�)'���)�4����D���U=R�}Y���tiu �sُ�
�C���ÎgVBӍ� L���u��O���FI���	���d��)q�lr���|�r�ۯ�^���ޥ�[7�d��j6̢� ��T��N�+9�%@�hKۏ�� .�k8>��D�5�nة��ko��O��b\��}��7/ôV����/�A+�QMK�x҃K6	��p戮\2���7��(}�<���on�"�p9�c+�E2��#9����=v �#�0�R��"uъv����c�&���{c�$/f���s2�W��3@^�U�Se6�����$����R/ܗ{Aw�0�vī��wp!��lv��mc¥��˔b��<��ى��ui�UȊi%��Bi5ۤIЭ�����;��3�e��n�c#oq�x,�S�|zӬͶ�{�pw�!!�d �O�eY�9yk\��S�b�š�?�����r_�%i0t�ksOŦ~��2+h�ii)�K��o�`JCvܖ����!�ո�{o>Z�_㮷C�� |b�;������%��Q���S�3�C�����O���d�]�pG�}J��6������VMʃ��*�c�71�n�;�v���9�N%����B���x74��f�"ʓ�>���_���p�.?����J�f"�g9�Ḭ/��5<d���Q�.��I<m���{�g�pR��Du�j�,ܱ��#Z|�cC�{u�R%s
��o�xr�������'�%��M�B'��T�W_���9{��3".�hA���0�"d^#~٦�� �2���u��O$���~���t��-n��`@�P��3��ݖS�5x*�~P���� �Y�E�Uu��^��w�F'����h)&��a�|�\*�f�A"ZBcs*��H�S O�ۘW�E�m{ħ���P1a6�4���7����5���,��T�l�3=M��{P���G	���J��v�{J�^F���mQt*3sB���Bd�%*j�3uNƋ�X��P��^~tGnF�y��>�P�����*�#�u}��|��j��ʹܵ��RIt��>�5�/�`7�Q�����0�N���\�Ƀ/��O�/ݦV��k�=���Vc����ܬ��ܼn]�zM��L�th��KO	#�U݅�6U���"ϝ��&��*��:ީ�(':��E�E������u�\�J�r,ٍ����+Gq�3`Ux���W{t�W}�%&�/q~���2!���������;[ȓ���
igiX�O �Hr�GU��.����nZ"�^G�U���y���'p��q����%�r���^��CJ�ɲe��)�א����f]uU(�ի����^�W�;�#�E���^��D��_h��&�$��ْGi�N����bXS��. ~�³Z:��\�h,�(K�i~��ѬB#/�A�{\�U�����u�l\��9NA��~S/!-�q���!K�Vʶ�qFBwv�ŵ3�UP��]J�}&~YSN8  5�M0^��li`�O�����:�7#q�؋�3��L�-�R���G M7�2�������/c�_�t��e~L5��:�cm,%^���7g�Y�&/�Ey� 1<o�Y�bld�����8x���
�|4��Dj�H ��e��7�
g�y-�GsKSQ��<�Be�S�Է����u���,���\��.�������r�TԿzp�`o��'��ժ�Ecc�\���������*��_�e�� �,`�夢f�I_�(Ѿ��W
����3���n�!f��tzh�O�?V.��<�8-��������\��;*�a��_A'�Ԡ�.�}'����Db[�u���ڿɶ����RP���u��U}f�aw����'y��`o�]wp�qy�.��)�-���'����b�m�z��H��q�Zoy�˜���~ʗ7Do���eF�U��_�������Xp���M�^Jk9}�9�2�YVP#���t��бb#kq�����j۩a ����g�sqC���4��)��Ebz�hzǺ'[�V뱧�.]R9V;�D�^����a��k�XH}����\�`0�iu��s9�m���J<�Ξ�I�����#|��t���S_��M�k�(P����\�y9�a���a*��г��vy%�	<�X�L^J�/�F�������O{�6S���UOi�����1?�SzڿIJ������� ��.��A��hF�|õs��Ɩ�*+�?�3��˻�a|m���P�L$*�SfFtp#��㯑�|��Arv�pV�܁A�ڗ�q������B��Td�l��W #O`�kX���;���6��D�j �|��j�ք�z���^���o���G�p&X��e��O��B��w��E���iC�2\��?�el � ��L����ڢc���ܮ��A�U��t���]\�H=�v)�	�c���u�]o�ċ�s�V_�Rh�`�.�b��޷x�)uެ�R�_�����Ȋ�z�۾\RJ]R>���X�i�w���5����.�Hvy��L_p�x���6����i�u�R�Ā啸����t��$�Hln��H��J��˥ݣl����y�g�F������R.V�DF�l" ��(�B^����Y���'�q��~�^I�Rv�^�uU�������7��,����Ӵ��>���S���1S� �E���R����I��ؽ�e�_���+l��k�iVļ�l�N������Bd:_�_�����μ-���� ���&���{*-ҥBĳ+��en��[M�kU�볺}�ټ˰C��U��FA�8E%1̦&ܙ�s��(h����Ƿ�Ȁ����Ӎ��=|)U~��*=���5�sw���%[�Ak��x���F*��y��0u9��e�&�	j�r�-q
I n������:*9���s�ZFɮ�#��!���d#~<�ΨG.��W�^��aW�������`)����ƌ�럇�1�UE֏�9"q�p�M�L��}*gn�2=�ʶ
�҆�O5Z~bjs�*Z6KtN���(�&��__���������W0{�;��:��|G�=E���	�.���)��Y�I"��W5�i��_U�W�)�@a{�3_y�@���_,c)�/���h�,
��S}88�LIɗ"�m��o��|/#�����t����'��U�Mh���@�}[j��y�n��A�Ĉ��W�����ʫV|m�}�[S���
g0�BXL��g�𺛩`����j:�q�}���Q0�ײV�^�*9<*�)��;�^�`������|B�x��b�(��8=�=
*�����e�]��sNK�ou�h:�!U0my=�gAG^p��r�����'�e��eÕ�y���q��>m_{���/����xi����/%iV<芯�yBd�o9��Vb�.�)"��/�����a-'�W?�ˇ�6p`e�W�cYCgPB�d�j>h6�pu3� �0�?�Ni'�a�e䌈��f����g�F��Al�j�S>��U�מ���Ѳ��CR�q���x�.|��<Ϡ��׊����4_��.�^.ҭ �h���a��6�W�
������Z��C&�w�(h�������&�4�ל1O�N]|�0�FHO����\�`"Ǌ��*����K]�K�?%��y�(��>�7��;�Z\��vsUi,�ZNl���	���G��2�d�-aщu���V�Mj~��\��H�j0�Gq\~��h=aȅ� �;$3�o2F#��2ɤF�D�0�3����G����Ud�����%�fp�1I�O+@q��c}'� }_�RTd��� �[7��F��؉{�d�M K����)��>��r�Y�=" ̡���ϋn[s�yvcfQY��?U�<����~��yR��O�$���<;�H���\ߴMZ�Y�������go�V]���z�o$�b���D;��-eP�?�8Z!: �E�^���"wo���L�!��C��'�1�?�Z �W؏����Mn���׳��6e�*����C���ON4ՋW�Kۦ^��]���)_��%ˈ��M�||�)�&�K��nH�W藙���S�Ut�8hh�[> _�d�Zk�(�pS!R��E<�9��;r�ĭQ>��cQ^=��(���������%r1�\`m�@/��������%�^�����:�p�P# ���d�3�Ǽ%w]�u�a��YH&d8>�ꊟ_4:F%�}�e��7��#;����
<�^����n���c��,�w�ZH���,�=�b� \�nZ����~��F�/�d[u�y��/p9�L"C5�+�
.
c�;��¬�q���ND\�y�		������X!q�/P���t�[�
T��B��sr�o��b[�YE�x�(�ʠ��Hco�:�<�gX�c[x@�O@wc�)��+�Q��Y�`�2��$A�S��1.��+�V��Ϋ�ԊH! �it�7���y?����"x�uU�h���ةE��{��pB���xdr���B�j6���D�ߍDv�# �{�R=7�����RB�9�D����=m��z�z�/��oC��aS\��U	�8YSK��?�G2&Kp�@�tOcjJ�A��������YJs�ĊO�i@��2�b�+�D=���:�jX����������AJ�B]�XwN?�[�����^��Iܬ�r/�[�PW$53�� ��Nt@M�������B1�[K����T��\��%��R���_���2]�Fv��\�Қ����΄����f�l���S/�����Xr���g����E���:�f�b�W�y��o@ ��� ��yBչ��߸V��ҽW?W& N��GK1Y���J��/��a��b����eO�H�=�|�`�����q�\���bF�Ѳ�Ŭqb�ƃ7#+�+�[�K���g\4?<3���.B��J4C�\���m7��z�y��l�s+�ш�Vuo�BH��Mz� {�y�\��/(�0$k�ޤ�ĔQ�Cʈ＿���%���  �.#�6_�Tw3=d���H� i�y��0/��4볩�	���s�E{e3�_F(^)l�
�e��@����g9��#�;���nBo�~�q���`I娶mٗ�Ŗ�f�=nxgu����_H\ �i�$+��H"\xӪl���VZ&�D����A����M�$��X��of��mv��o`!�Z=����v7i�~�ѣCI�Xa�x�;�'� ������]mi��$P��ج��*7*� (1]�P���V®8�z��@O�b4�T+;�o�p2�����f�1�����o+2{����g���T(.mr���X�^Lٍ~�e�5~�c�.
��"ǁ4��߁�A��p��?7z�Ѫ�V7�[�K�f�z|�#�L�k��@�?�iq�����:�b������՘��]�-���M��~;)�e�V�D�v�i�>%`\3̧|L&�O�Wd1���v���3}����8/_|��&��R ��H-�0�����nP���4����:��ԩ���K��ls\�f�fl���=�p+�X;��/2��ÿ%/���U3��� ��c�u�l��'!�(-C��|Y�����`ഃ���P��>� ����A��/PK�0�9�  P  PK  ў,J               226.pŔ{4�y�y'�	aBB��L%U�F=�#�Gu�t̔����]�,ZT���c�j&f�������JT��iI�sb3���������s�~��{���Ͻ����d�����  h� �Q�@��8�@ P(��VYIQQIKM]K���!h��Ds2Q?	��X�?`aii�K����6�YR�.�P(%E%��2���ף��!{`� '����u ��}�@o�-@`G Q
��w� ���
�ͦ��(��g�Wg� �c�Դ�J$ɥ�M����-46���NK�ЈL16��:hmc{������I_?��S����~�ɧ�"�>�O`&^H���̬�va���k�Kn�r�������Vݷ���nc������NAWwϏ�C�OF����ɩ�3�s���׫o��76����@ �{�K/̮
�@{^ 0s� ��Y�՜��u}j�RP�І"�N�h��(hXNJ��ޚ�{b����?���%� ���A0�#�RG������C��6���z�W1�J����VcYbp�˂�JX�� g���Φ|}�æ  �n�/y�&;�w>#����L��V�cuB�("#�$�^�p�����s�ǖ��H���ab�:���(�9���W��(Z=כl�u�j<����cXHe�e rZ���Ϗ��gyƄ��`�Dy�%ԎҖz+C\�G�;��6F����Mؔ!��c�<ot��E�?�8�x�R�r�e�y$��i�0)�(t�XY��nI�2�^�q�:��n;ޝ��t���x������b�Jٔ�h�4�ٸ�lj�r�8�͚Y��;q!�?�|hc��]���э��/)�����|1�a�(�Ty*W�OZ��Y��CD���V�p�M!c�4�c�<ҏ�a��hA�C�0g)��)
N\�.��Z�as�ٔ
�T�	���L3a��.��Sd~��Z�l����y��{]�7<�{ftY�+4�y��C��i ��r\���Z�(��$�w]Y7���Վi���$�:~�:Ҝ��&�8��f���6I.>�L������B����H�D��{��o�XYxR���hS���G�:�:�y�ch#�ɌD�,9Az;�{��1�&�٥�sw�����s%ه;���qU?i�y�V�A��aݧ]�\�Y�^��s����<����e%��ލ��H�P�E�<��]��k<��Mw�#E��/L'Ue��>	��m����� �p,n��4��Cr� ���a��9�}BD�;�Oo-��s��m��o-t�K�N���T���ҥԮeInx�5��)�g�vۿ|�s>^�$܍?��.����������I��^����R�S�ht��W�͡f�|>A�4c��pe�¹��A�b�3O;�V�_�� X� �-J ��O���������t/*��B��h�<b:�d}�'���d��|x��u�x������a��2���������h���芴�dP�������r�����P�
�'�|�/c0�,5��%�{�TM8�Q�,͹���ˠ�z�����6p������;�SPڂ��a��O§:��ȕW$Ϝ<��M���;�i����g+����T�.�^�Z��;	�lL(�ڐw��G���k�]ꤻ3��r��T]�&t��KJ4��sD
�K�2,Zj�,����ʄ�RSC�(��!/e��'��Ꞟ�{�>��7��_PK\G�.�  �	  PK  ў,J               226.vec��Q��=��k�؂-�b+�b+؂-؊�؊�؊���ݭ?���qɰ���9g"�|d�J���N9�S��)�J�*[W�*ըNjR�کu�.��O҈�4�)�hNZҊִ�J����=�H':Ӆ�ޥ�v�=�Eo�З~Y�u �`�0����YY�Б�b4c�8�3��Lb2S��4�3��̲G�us��|��E�B,�%,e�Y�Jb��b��5��u�gS>6�f���mlg;�ef��a/���r��f��Q�q����9c欞�G����e�p5���׹�Mnq;���垙����C�'<��<��0���+�׼�-�x�>�X��חb�����O�=W���gi!~�o���� PK�YErj  �  PK  ў,J               227.pŔiPSY����$$����U"(B��ЀQA�i%�`I���n	B�D@0��DV��Md�6I����
h�%�M��g��4�LM�|��_��=�s�S�j�j?��`go�  ���Q(���0����qX%%����M�-Zĭ[�m}Cm�z�|�S3
�B4�o�����n
y�' ��*a5p8�A���j5�� � P@���*�Z�}*����@�T@��h��|� B	)( ���0�:�TUP�1��6Ӽ`]�!HW�;XT���2�����|񥆦��6C�v#ʞ����[:lkw䨽�	���n�觙�>�����R`;�r'�Zt̟by���)�7oݾ#|�����������I����ں�"����6ɛ���]���GF?��OM��f���ּ@ �^��KU�@"!$��"��6�"t�PjT��ڬK�P��ՠ�v;O�3Z0_�S�L��}6���"�+���ӫ�B�<<H�&���#��4��\\,��[4�w�Vԯ"�J����x��%�3=�(c(a��~ϰB�u���B>
O�~� NgY�U���+��8D�'_?2��:Pu\�'�27�7�~��}du�(q4��ӽ�+�C��"� �.Uںy�z����f
,^F�|�`�9�[����%�4��J�x�R[�ZBT�������=�<�]�.sX ִ�2�4�_�՚�]����ǌ������~.�4�}\?�Sg(�կ�;\�0Gu6�����~=��Nۚv�S�s]1�41�{{G$��p=ڕ���K�G�Pm�N�:�́{ΖM5Fy:f�1+;��ȭ�����h�3#;��l�E��V|Q羑[-�>����v9r;�Y�N��i����w�u#6�9�1����,�G�mב,�ڊ���=��Yd�}y���&䓀u��D�A��O���{��H%W�@bq3%�Q��36O%��7=}G��K��\8]K�6��#�\����2]r�����5'n�9�u�/�/0/�;�Y�K��~9�6�\�|Bɕ��V���{��7�2����jn\����c�������ɮը�2����_p��q,+NK�%���z>G��^mS�-�|�tކ�f�5sP�Y�E=��T�5��A\y�v�q���,�
+y'^�D�z�3y����@O�\%A|sv�lO�O�. ���P+���uk��><�F��'�����:d{��_5�]����FHV�hk��/����n���\Jړ�����Y3��q.�=w8���c,�h6�B󜈦���o9;�l�jz�Tk��cIB>�2ݾXR��߷e�}f�[��\a�	�9�m}�=�4�e��ἀj,>���g-�#�I����W#%|��1Z�i�C~�g7��$D���
�:�nKn��ҝ���b�h6GOD9��,ˏ���I��WN6N����C��X_����,Ӎn���R}Os{�[�H��R怨����X���s��jD�8�onl���i��(��wT@?�uh�
+��T���U��9�g>c3��4��x�(�&1M?��9�C!�ۜ,� ���)�^ZW�,>T��w)I4�5�޲�������P�G���q�s��m9�S���=�ʜؑ>t���k���S����s�z"��a����/����ӛQ���-KRm"s�����b��2�eAI������K�ވ�-���eߤg�r�6�?�O��οPK�K��  �	  PK  ў,J               227.vec҇�Na���y�絷le�&�l�)[��&�l��&�����Q������sw�v:�Ӊ��"s�PJ��w�Q�
TLYT���\��T�:5�I-j�<�h]�Q�4��iBS�ќ���i�e�V�ўt���B׬ݴ;=�I/zӇ����:��b0C�0�g��#�h�0�q�g��d�0�iLg3��g1[�0�y������,��X�KX�2��"��J]�j�5��u�gm6�f���mlg;�e�[���}�� 9�a�#z�c~�q=�INy��z�欞�<��%.s��)�5��nr�۩w�.�l��f8?��y�Ӓb<�缰{i���5ox�;��|�[��%)���[!�w~D���y����I�?PK��@�e  �  PK  ў,J               228.p��y8����$��!�P��hp�PT��Ш^b�Vq5m)7:���jKCE��jI;el��i��c��EZ[���ɠ21ϝ���ֽ���}����=�9��9�9�q���֚d�  �OV����������.*�@I ���R�_�����1:ʪZj��أ�ZGt�x����q#=S}���" G�#�h=y����] R4
��* A�P$�(	r
����!P����(\L\0�q �P*$�	�Q�> C
I��ZK��ET�(=�HTͲ�{���F�'�:\L� ZVV�0��𨑱��	���I�����׳��(����x��կBBî�w#>!1)��~�o�Y�9��{�%ߔ��W���������G�{�O��}��Ǒ�F��'&g�8/^�/,.-�}�~}�����@���_z!^
��!a��0!]a)��7UZU�&��d�u��������`����f��]�������$����˃"�V�e�]�c!�#$*[L+ɲ3�ͼ�AH���+�V�ʝR�H�*޽����R5�����ѱ,Z<�l.�	B[����T�A/�n�����"�-�=�f�4���&I����#ـ��1��Ď����v0�f�W�}���)��,�.w�i�/�b+�R�G54�ƫ��MW�ЇK��	Y� C�V�#Q�' 'x���#g�`ŤؿKgR>�X��G}���õ���j�]4��L����k�x���#��d��^�,��xt177N�"#m�~Y��6���$�J�鶵�~U����1��*Yڷ�a*����d�}�a�|�6���1���H^�]m�[�xt0��v\z\�>k�gd�$R5�+8�
�^�x�>j��p�y�b����F���J������Z������Kc����\�tU���;���y���9}��B��D�s��e���oMa�8z`�+���rO�/��2�.��ҙ��j=�6Ԥ~�K��-�_�b	j;���CSQ�����upLv�����m��b˾���F�|`�dP[o�<��tV\W|Q�j������E��s��x�p+>�E�>�^�˷��˗���ڑ$;���8$m�ᗼ��Ev�vÙ/x��F���TӫG�-!��5���#)T
�MU�$��i�050���?6�7�����+�Aòb?�`���*���iǞ(=����嶄GW����ή�H7���}�J��d#l׬��m���+UU�,0���)�n-�sV��A�_f��9v<Z�U��$fn�f��5&���3\�����^�Y����م��\,[0�Ov���_~��n9�����7v�����_ɑ<bTk�r�0��+k~��k�l�c3o̭5k?�
_��Y&�v�vX]lO�)�Ԉk��O%�!Tn���M|��j�b�����c9�4�͎q'�6����V/���L+jg��l��v�;���r�Dݽ���1r�����S�K��9��i��,�]��������:|ʌn�i�VƆs��A�۴V3����9��V�-[����DZ&:S�:|��O� ;t)7)��I���2W���U�,�B�y&v#w֜2���x�
E'ϐ�R�}�+S_3D��!���epyS(�|�Ɯ�yT4���'5%OE��&��� ����g��ikQI��1ʬ}��<aIՏ�����p74��36j
���	��:�6�����G?��z��,��|��X��0��^��w�pb��+J,�����$>�X�X{��Ѝ(�>3J�
0�c� ��ʟ�PK�*  �	  PK  ў,J               228.vec҇�Mq���y����l�d�M6e+[�d�M6�d�M��{�Q����tz��u�t�NDV��UF�<��T�"�����bWչթAMjQ�:�MŨ��i@Cј&4��iAKZњ6��]�E{�@G:љ.t�ݳ\�О��7}�K?�3�s� 3��c8#��b��fc�x&0�ILf
S��tf0�Y�fN1��:��,�E�"��X�����`%�R!V��ڬ��l`#��l�E�����`'��������� �8�������'��9�Y�ٜ�\,dqI/s��\�zJqCor�����n��=�������<�)�R.��^���������|�#���Y_���~�{!ŏ|����W���S�PK�"g  �  PK  ў,J               229.p��wT�Y��/=� ��H��@��C��BpGE�DYF��.�iQA�"D@�F�"�08�t���U�2@(��F�ݳg�;���;��߻�>I�dPp8p�  B  �.@"h 
�@"�($�F�d0x9��,����ūo'i�oWSۡc��C�@[M�l�o`lbffFҳ����545�n�h4FC��#P5�4��qH�8�ȁ�Z Bq�� I�	?�� !P�D�ed�� �B`P8�f��y ��+j�|�Pby!�����[�(m�'/�]�guL�s�2�T��;���3�=�V�4:��A�!�c�s=��~������+���!�a�#"/�\���OH��)�vjڝ�Lރ�����E�J�~WV^QYU]�������[^wtvu������GF��'&��?��/,����"��(���U/���Aa�M/rqs�4A(~�Bz)iQ�Qx�[�O^��M]f����l�1�~�T�h���8��ٿ����`���yP`�>"�9\r�����e-P��j��!jnf$�60�]S���ߞ:������fݣ�=hr�u[�Oe��x*C�]�6r��>������ �*���R�ѹ�ό�Նg�pC�3�j�V���?�A�1+=����k�{(b���_]�����0is�w��T��Rl�潃N���>��Q�.?��L�@L����ލgg�x��}ˉ���&*�2�w}��z�����Dĭ��Fپ������7���-�T1�\�#��T�X�MDSx�턋c^�O-��.kR�"x�x)�� GQ�7�x���v(חn�B��s�\<ȼ­�#_�H
��]=̏oA���+d�D��@D�s��{y�S�`����,h����8V��l;C����lb]�d�*�˝�K �p�oT'u�/g\�]`�e���h���)��è9�P���Ewx�"�K�|�0�*�k]>�+t"R[XU����Z���
�*����x)��1��SI��Y��=��?�>�&��ս\��Ѿ�εz
C�R�o�^Ef�_,!�H���3K�	��	�>��D�ׯO4��­l��f1Lb���O�zJ��[|dO}l�z����{Q����(ApPN.Z��Hm��bʾ7=���6�J���m�S(�6�rϽ�L��Ta���]eO��Pi��IN`��n�D���*[<�ы�w?�m𹱮wG��#�*��~w�,�C<���j�9��^�t�E���X��P(��W�6O���3�z�74�����m�u�He�0�AU.����������HK�QpF�C��ZM�I���}��?-~����X��bS�[�j	X,�yU������y���\�)�3?P?�9h��=�,�� �r����=�	�]�}@N�u	�
J �!���8�=��dg�M~�H�������s��\d���nh׵�伹�@�Ϻ��ڍr�cM�	�h����vK킐��z�)m��QjTP۴�S?~�E:ׄ��:'�׼��o3�0UM��؃�MVOg`M,ȗ��$���I~R��_s�6�&z�~������*��1ZE冬�S|���y\J�V�Þ,�=<ς����!��}�����,�u��A�����xq��l	�fw�ex(`��O�3ªMe�0�Ro�G�&�i�E}�ݜxng`���	�i��|.=@��g����kY�ۺF��S�_R:�6}���;�
j�1Y�C�=���P�6�SG�+E�1���'y��[��/d������Dľ��Ŷ�·�!Jׯ�Bn�Чs�Q"�8�@ӵi1�S^zk����E��7PK$H  �	  PK  ў,J               229.vec҇�Na���|���[��e�M6ٔ�le�M6�d�M6�{��G���q�t�{:��9��#s�PJ��g*P�JTNYT1WպթAMjQ�:�My���4�!�hL�Ҍ洠%�hM��.ˢ�v�#��L�ҍ�YI�О��7}�K?�3�>u��P�1����b��fc�x&x#u���T�1����Y�fN1W�1�,d�Y��T����dU*�j]�Z3�t=��&6�blѭlc;;��.v���^��~p�C�G�����'��9�YΙ9���_��\�*׸�R�Л��"n���qO�{7�<�~�c��g<�/���������|�#��l�/%��U���G!��H��=����PK׷%�h  �  PK  ў,J               230.i��g4�Q���c0�5F��n�A��2��ѣ� b��6ZD�eBD����{����E��]�|�����i�u���}�.W�W��M-u�: " ���f� ))�������QP2PQ޸A�BGO���
�`gec�����}���M@F𮨘��$�_V&�pOBR�?�����)oP2SQ1�s�q��?�U@KR�� n���]}���$�� �C@D`bR9ōk��� &"��_k__�bZ:.1Rzk�'�xHR>�jm;���.���W(9�-fV�;��B�R�20Y���54ZF�HS��([;{�g�N��/||_����GDFE��&��b��32�

��KJ��+>�}�����������ή��ѱ�ɩ�3���W�����7����O������A�S��\��\D��`b��@D/�c@KL�%FJ�b ����!cPMʯm'�0�e���`��ͷ���&����"�_`��k�����������}���վ0l��LF��,��,�@����9m�O�:��g'y��Z���<KT&��/y���C0�V�B8����Om<���F�|N���bfo+���ʚ�E��;V�Pok��r���w�_L 4	����[�m����9Vn�	�s2m�a�}�h.�ﰡ�t_���u�)N�x��	_3*hn�tvID&�Wr@���w�K���Dr��Mq"��V�xVn���·f@��_�ߪ�&���v�tp �K	�	��#�_'����z-6����۲f���`����������wesZ����/��/֫�r=��-i�~M�cO%�w�/t8z=�4�ICUe�L=sqE���)�������~��EZI]�u�1��1�G��q�����^[��3ZK��*��W������8�j��i"���ez���ok3;�P&�x9��g�zS&ɒ&�������E���?�7�#Bs���j?�7�KR�K�g�3w|�
�Zm���V���k�B���S^uߐ�+ �V���⢪�w��K]���D���ika��nFs�����Q���nuG1Pù���j�G�7lz���ܓy��|eb�����\�/&d�;�1�Cև���������2U,�M"7���B�|U-�}�|����Xd[�7+�w�y���.9�m�={4�Q��^���=a@�#}�w���Z�b�u����~f�~�B#�������]�ƠȄ�Tm7��b�?zl繻�.t	��K��*�Oq[�
m�r<��O)Ryc���M�����(
Q��+p�`������eX�ĬT5�%�6W�м�8�=5��8�v�ʬF�ؗ�x��3��h�b���;��Ѻ�[�l.�%�o�|cxE�|�4}#>�����՛ge*8c<�yi�rG�ܶ2�������]}�������M8
�O�̝�{�qK.�^;i�)w?끿��q�w�Y��رݵ�eͤ:�^�y��^�s�NY�^��g�z�Yۺ�Qg���_��a.:�c7��&��G?*�9�@x.�զͣ�à�r��^C�ƈ����H"爝��}U���[�d0�6a�VE-a�,�qN21�FbA�)�]X)Ԋx(�Xs��V�h��n|������=r\6�ҡL:�-\L�ޑ����M��jK��_H�澳�W
��f��il?��ɟ���w��6�˧�8r^pd��~�9g�sc9�3X�2yTm>L�b����U_T���䰂E�"fv�Y�v�ӄ�:�YSס���0�(�w�Յi]V�QUrIѵ�z�l{8����u���4���M]�̑o�3v���M
�,M���[PѮ��'枊��D���ǧD��Xa��l��KY��Պ�-�K�&˩��S�ڧi�4���%m��N�ؐ����/ {�����I�6ź*��<b.���Sn빲�ΐ)�Q�r��\�eJ�l�3)�ݥ;�hqɑ/������Sr)x7�%YO�cH��Q�G��`<%�gN.!���Q=I��r�1�O��OtBY���Ë^��qڃ4�Z�T�E��[8�VOP&Ɏ;���=�w�r�D؃��SnKj���I�1�_bfӸ�O8��*�ӍG��tu�G��$)b^Q��fQ��4�k��['�9O�ve,��;[DUێIy#o8�2{�VwG����߸ �!'�W�S?)�i�5T+��6ϐ�����1vl�q�09�ЯGZrw{�)4��W�K�Ug3��仞���0�B�1�����*�0x�c\�d�풀{�������~ ��� �c�.�vZ(�ן3�h�!]��s���qtzG���|��9�4����'@�M�Sx1�´r��N�f��>�lM�WM}[$3��m��+f���Y"�X�"D�-���p��F�R�yy:���D~o]�U�_٢Gr����ߖSu�t��V!�%+�	7�qO.��xS����}tt�'��vC�Ϊ��"Ҟr�2C%���_:Io�d�:Nϩ9���q�K�'���ȭU.n\����v�X���k�Nx���tl�RV�Se�aR$&�k�ye�>�������G�x)�{)�*3�g��j��bq��7�>�NI16P*}�vO��h&I���7��n�"������`��a������"��I$B;F�"Y� 7u�8�b7���ŀ�Fy�ͤVj������������"8�Lm�j:�t�8&���C(�
g��>f�.�`�E���^��n�|J��9��HK��1�-f��m�&�6��w�F���0ơ�_
+����j%8qz���?��s�Xy��N�O낐9�+:7V�7�,W ��d$��}]����w�\��q�
]g�����֏=7�t.U@v����\�˾0Ff��y��Z��=<^w��K�m�E�Cf2�e,���e˚�S�Plz�����c[�5=},o=:���<B\�^3���Kp��ru����ߐ�d�c�;Ů �mT�ˤ ���5^O�ˁ�X�D��ů�u�21�;6J��u��o��iȂ���
@��X�l���e��[� �ըzXS�]��e��P�/�cm'���;��\5�'���ӯ���<�7"ߛ��hK�������j��{k��S�#+r���Bh��*�COU��M�|v�{Dgjii��v�-��i��P�b��0���#Wg�	y��{D��N'�,>E�����>�8�P��|ó��!c��Ch�&cz�sv��4�ƚs��c}�2�Ȧ�cW;��23��⇽H�_�c�o��k`qu�aeN�'�_!bQ�0�Q㚶h���1�)�g�r)d!��E�+lK���	�ɤ�5�y�;UϷ�?7�y���]�%�z��3��� �Y���!|�R�R���i��Y1Q���f�2sʯ�KK���@/S�yGS��J�繜�v�b��Up��\��."t|UQu&4)۱�/�ď�]���U���y{1,�f�;ݱڝ!W��:7V�~�֕��*��n1?ep]9V�Y7��U�r�Kd�I�&����Kr���ݤ�l��E��R��^KB�&.y~p$wJ*��f��HS+��'5P����r��]S~�hL�)�d�(��β�T� ��B�C��Z���5%f\�B���=s2�6�[0�ꞝz�վȭ�G�3����+R6u²��*Iw��ǣj6�h��A.����%
�x��U���c׷Z�~W&"�ަ�B�WY���&s���N;��	?�pE�c�������/1p�ة��R�_����|��L�.������ѹ���Y ���lr��x�Ǌ�)l�13��9�#�َX����o�vF���o��f�>:��l
�饄R?�r;-���O�}�^NF�	����1���,3�H�^)��uA�%��q��E���?.��-y"�5
F>O�S���8��|U�7�pc��į�޿ʐ�����Gb��C���yNk	��z�n4<�_�r��v:H�0;d4�ݶ�@�E�aR�����d6`RI9��1*�ʿ���g�-i'7aR���Lڡ��|�M٩�����)�����T3�cw��׍�:��e���C�?�H-��&��A�{�+�l�K�Ğ�N)JN��e���u>�Q\�=�{������̿��,�^�����ќ�T�k�'3�`x��.��"���}{l���)L�%�ܜ���I��c2�m��&�7A
���Us2��wʓjV�Tȟ$�;%�{Ho�Ѩ?�P�<~G��
�:TxF��pz�7iN���>�*}�;�VDc-'Ӥ�0D�}���~:A~��}l+��@;+��ۿ<�T�U��(*ɓ0(��@$KF��n6�됻S��]"����v��7��u����k�QyiK攥��b�/��7�s,�~�"4��HQE,e�)_��RӍ����f1Kh�ޝ�2����)�!�ɦʱ�<��.t"+l���V���s���c�+@���AA�����;���f�u��/�5^�1%����S��dά�jKg�{�>�ٕZ+P����"Z�xMG���`lѡ�х���;T�Y3*�����������ԟ�s���O
��1C�c{7�7�[��s���H��"�խ8�_���&l��d��.��c���TcCK0��UxR��9��Ǎ߲媥��$q��U�g�֌����ɔ�kB����]v�����w#�[��LUY���[�o�T:^��:LE�����}����a���N�2~fWɀ#4���4�*w�v�:�U2��0���fv�[LQ�:o�<���gy�r���[z���Ȝy�����i����u���7X�M��v�e��i���=��X���:���˾J-��{�Kr�_hP��r!F�����9�9���5>��7�~�5=�{��z��9�dNy�1�tViޢ���S�9������nC���!���O����
���0�������0������~~�@��=4h�,�����pq��8L�P�ȸ��Uń�M����͆�Q>Ŵ����ɹ[Z�Ί������ǋ���\���)�
Ɔe�)�	��m����mxY���D�%��o.Ń!�9�M�kWI�+:d�x��ՎZ�EgCo���UivюY1�Ky����WT͊C����	�r�$V��UػԙNӼJ�g=M({�+KW��������M2�g�-���D��v�K��qzۚ�y/��7u��}ąM~zX�����o˛8��Ѵ�x��Q~�G�6��gSR:����koĳ�#�;Gt��[?� �j|0�F��O��u+���*-S���+_�;!��;����L�#4^/�(6v]��j�פ!S��<h���NM
�m코�)�ֳ����#t�}�X��J͞I%���3�i�*e?p���M�x<��oaJ��Ⱥ�
�RL<��]�b�g�v��3ֱw��أ���w�4vCɆ6[tӽ��D�+���I�Fc��C�l{[���YƯ덡p�Ę��0Y`W#`㐅���-��f^ƕ���w�~i�H\�[�d�g&ϗ�@ɇ�9������o�堶�V�믑|� ��ѵ@ȋ���u�n�����p��9ߚNYg-��R��Ò�t�p5|�!�~p��P3����%�9���l��Ky���>J�=�LY��9yJS^��uh�ÿ�����!�Y�u��T�
��ػn��N]��ȵ�Ȇ9�uT�m7pI�u���~(aKK,�H�˪)�
���I56^�o�õ7�shF��4�$糊ʜ}o��9�5-]���o�3�T�c�h���/Y�k��J���|-�
�eKH��L����uI8�=����t�"�e�w���Q!E7��ķR�NCB�����7%e }G� |���DVW�?�a~^,I�(`��ӗtr�,eQ������A�_�%�Nw���DՈtI�#��ժ�ɝ�gcN/@'�뗏�s�4��Le�'�G�_�������
���
�]�������D!��!XA�q�2_�����oI��������΋N�+R<���ipmb�T�I\E��>�D������d�~��$���5O���5䔟�T_D����!��!�����]
�-5n���]�:�5�/s<A�^|q8�pڍ��X�@�0�z1�Q��"��ƒ���o���U��Px�� �H���1���^�.��	��Q��`�+l29�y�i��	�4R�Ϯ�k~+]I���Msp����^`�RT!E��L���N=W�L�v=��~��/�p���1
�6K-8f����yho�T�����p:��F8�q��c�׉�<���F9�r�?z�?��,u��A��-�P��)�d�i���hQ'���T��e����S �sF�L����i�E��)+��@woA�����6b�u:��}�<��j(G-����b��{^�A>��yx�3�J���f�!D��V�����\q�]��"!;jj�D��X����������������Iʔ��ѣ��a��g4�/���_&�0x���hV?�®�1�N�p)i0�f��	:G3<��+���*�J���z0E��|����%Rj�ڿ���u�RR��^�ܻr�����;������}�+ xJ�b��K�m��m�99�i�ԝ��j��m�4q+��9�e�_��h�:DM�}x1��
�&��;�9��hn#��&��<vs�n7�q׮2�P1�a�4[�
	���ƒh�J�4nŽFlԲp!x��d�O���{�Ip���[�c�7�^/S.FK�V�?Pc0�37N����yϓRtƏN5v
�[W��0�GV�u�:������@�ph�m�kG�Q���jnbL��cQ��:���<?L�%z��Aeygj{���?Q5�v
�yo�^V��O:�`��$\Ƒ_��>c��q<|V<����j~m�T�Jk��h�
*�m<w[/S!4?Ҁvr���Ni?�'���¨wA��U7�ɩ�d�سf�D�!`F*�~����g���m�	�yh��G<[H�d|>�����ɍ�zs2�4UMUw��4U
u��Ъ�Hpl�~#��G���M�n<��Jr�Y$0߮A��~���#^��<o�Ő��vtG'�6(j�(1�FOM
b�fו!֚��Nz*ej�np��SW��P�V��+�5��o�~%5Λ��i#T���]���$��cR[p�
�
�W�H!���|���@+`��&������ټ�0����]�~�LlN2jH��������c���h��J�0Q��f�2����O�L6Pת�9��%�η/��kq�_wgG�8:�(����f���	�ļĪٌh`1��x��r7M�Y�i��cj8�%�b¡�m�K{{�rb���H��s=H�f�*���E��q�������:T��� e�Ñ9a�� �b�;W?�PK���D  �  PK  ў,J               231.p��wX�W�!"�bVkM �0KJCP��H�L*A�0D; �(C��Ȩ�Bj�"��
�`�XAV���ނ������׹�y���W< ��l� � �$� �à8�D"�Q�m(���
�1�*j;UU�Xu�=:���X,�Hw�^�������Acҁ=���" $��A)oۦL�aq��9� 2�� < ��� q�&9'�1�H
������dC� �� `(�dY�< AC�qDs��$Oǐ87�FE��9M}_F"RZ�3��U��u�����Z�XY���9��us?����t�������"��c�������vFfV�՜k׿��,�u���������5�uM�-OZ��킞�g}����c�����z�zz~A�����K�7�@ ����\h	���7�@R��(��7��O��Ƃs�׈��w�S�etK+i�i�o�}$�4������`��P`�dx`4@�J��D6!_�o�l���(ﴻ�vg��	��Yc��{�ǗW�� g3�°��p� w�����I�(���t�Kf:W��.��c�m�{,~Yw4̦uVh���o K|�ri�J�8+�(�/.%}1ڇ"κ� ޙ����4Բ2��?��6�Jx�r�-jVad�e7��q��@�O�<\M-I_��Ka�LX�K�;q�f�,��d�5�`��=��c�˓Z")�������+l���������϶1t�}�c���C�ꔢ����f��r,9ϰ�}����8tT�� p��f�yH9�_o��s)�iaX~P���$�|�?Q!����(�C�mC�.����=ܢ-����.�h$�J�&zNe���D�H|TZ6O�}!���pin�]D��}���l��iI��#h��ƭ/�*_#} ^�v��}xo��1�'z^���|�U	N�ͭu�pRMtʩ��3)�O04s�-��� ;Ter޲���z�\��u1��~�7���.�»���7��G�O;��Cs5���Rle���1�֢�+�Q��!zoqY��=Tԉ;eJO-���'w�a����`����3�rg})[ٰtܒQw����P�9F^��̭��e�ZF���mL���=���+ܤ
n�U�s�A���Gh�h�^�S�&��a�5ս�C����|�3�����;_�	�kM[����%�x�S�9�T�U���d�����M����+OâC�G���_t�sw 3�)�V|kح���oå!9t�J˴|eDn?��O���gf�Ɵ��3�H��پ�B�="���&��ؼWF��B��E�n/�7񮲬l^a�p��m��j'.��Qu�w���zBѸ����Zt���ް�s�{�״8�B�ꁓQ��p./��g�����:>�}�	Z�	̒#�V��a�<P9v@D�
��D-��y��@"��sA�p�Rq��㒽������������鎊�rǝ�&�C]���W�ƪ �j�;we�R���o��C��d=��i{�|���\�`�����boX7K׺�{�!ﮅ9o3�����UH��24��~�.ZF�#	�Sq5d�Vͯ��<L����ǰb���eÈߔ���T�ѬS�_t����tg�]�0��B���8�uŁ���Z�#d"��~����"�6�]O�cq�Ax鈎g�������qY�ե[}�����
���m&T����<�L��{�/�Y��C��w�n��r��W��5cP0��������T
�eK����PK���  �	  PK  ў,J               231.vec��Q��o�uu�.і�D':�z�Kt���D':щN��{�Q�{�#�'���˜3��H
��r���;��BU�eIT7Wú&��M	u�K=�Ӏ�4�1MhJ3�ӂ���5���-�\��t���BW��=I������C_�џf� 3��c�7�#��(�Q�fc�x&0�ILf
S��tf0�Y�N�1G�2���X��\,��,I�X��X�
V�*+�j]���4��z6��Ml6�E�����`'���3{u�9�Aq�#5sL�s"I㤞�4g�������.������U����eq��&�����Ҹ��y`�>�1Ox�3��Ŋx�zm�����=��'>;��\1�z�7���Y��W�<~��f�?PK��Nl  �  PK  ў,J               232.p��{8����\�DC��[�Z�aq��h�nYz�T��K��nm�2ea;;�j	�R��)v�-.G#�#�V-V&ոUk�g;�3�9Ͼ����}���~���}7G7꾞>�  P9��1�PA ��
�D�T�X�*����ح����GO�@0 Z�Y${s˃�
E���Ł|�ʆB��D�PXV[UU�lH0$�ϱ��T@7�
Ł�����p�m �����

�Q.�F��P(��a0��%�< ��5������H#��ŭR1v�s_�d�h���Bk��ޫcbjF2�G���wpt�x������p,0(8$�q*�tT���Ĥ��)^H�|��s�Z.�����e��oV����}����o��wtvu�zz������Ȩ��䓧S��d3�s�K/�+�k�[^  ���SzA`0(��BR��`pCk���<��mD�R��s���G�]�O�����I���[��N,��2��ؿ�X(��<(pkI���9�Jȟ�����|Ɂ�)��#�i��!�r�髋��~�\��dn�dlr�� GS=Uk٩���ǘL�Ѽ�wO[jv�ж�NN+��Y�R�9�~U����ݍ�u}�Q����,S�<��� ���D��ͮ%O-��1j<�eR͈�:���S|	%p�!��Cje����I�Wr�����zѻwJ��e�9!�"`�G�\�c�2���5���cTe��m!�,��t�Yl��xdU��k��ƼB(�W�As�u�9�EY�B��늚�F}*�'���G�m@F>�c�x���
�D�w����'ǋ��t�^o���ć�"
��=�S��j
�q���<N%�������G)2kױ��ef|/8(|�p5ob��@�a�_�axXɄẀ��dg��;�㐀m����6kB�,bx$/j-xR[�`��u*8�i�#�vs�h�@����ϔ��2��t�N�@�p�gb w��/7�'�_[3�/==^�ϴk�{��kF���)v��i.I��Nl�;��KaD��+s-���S#�jJD{#��0���EF�U�փ+&��u�k��O�Y��K�Y��t7���n��(fh쪥�%�;[%w�f̏6D�	�k�%�B��$�:���{h��Q"=� =�{���Sb�"u�$�q8��q� C �`����ɫ������;zA_N�Ah%��h�緲$��-W߅d��`d��v�s7s�������+�3<O�ۑ���/��Hq�[K2.*3=B|�����F�@�i������Ϟ�W]@kC���Ame�;��x�⯶:�S��
 ��4̡J��V_	�*oB��_x����
E�Hس	��-��
��-���_^���6T�Ms�W�x�_�N��$���#�#�ا��4Q�����H�S��E�G��V.�g��o��x�me��W,gZ��}ڍ���O/��5�P��Zm:l8=B���!xbQG]�����n��OyK�.�J�ںe�neTLs��"��G�Ke���6ћw�'��6�Ak`��r�މ�8����=�}���1w�{������E���v(���b�6�t�u���8��1�YyC�|L�di���Լ����Ū��?=m���#r���x�Ow��E�I���u3w�
N�X�
���c�U����ُ���웖�����[�Kd�_�����FX;����tf���6F^�lN�i�Ԑ&����>�?�R��Zm������u�r����_/���[[�L���2�a�d-I�S��l�M�PK�'�*  �	  PK  ў,J               232.vec��Q��3�Z�E�K��щNtb�b]���D':щNt���ۏ��v<2y��LNnH
#��(���T�5��%Q�\�ԣ>E4�!�hL�ڭ�6�-iEk�Жv�����1�E'�L�ҍ���'��$zk�ҏ�` ��Dѡc8#�(F3&�G����r�1�	T0�ILf
S��tf0�Y�N+c��e���.���b��i,�e,g+Y��j]��|�t=��&6�٢[��vv��]�f������� �8���9��9��qROq�3��\q^/p�=.�e�p�k\ϲ��7��m�pמ��>�<�G<�	Oy�s^�*�����ox�;��|�s�U�W{~�{d��*������Y�PKg6�g  �  PK  ў,J               233.p��{8����c.X��`��̸L�u1J���bHT�rI5��\r�ܦ:.!u,vBjkB�5ƐK���[��XB����=��e�<��}�}�����ޟ�W�� R�,�- �� �A�@���Ea8�D"P�h	q11q�]�h%����SU۫�J�C��HF�����dM������d��G@$).&./!!������t	^���	 D�J��"��Z��
�@E`�p%&�P*@@("��DD��pa������Ew�.�	�h�)�!����d�����(���V]C��[�l��Șbbq�jiu����)��N�g�zxz]��t���@Fе��И��q�	��Իi��2�?`=��/xT��Iɋ���WTV�7p�M�oZ�{z����?0:6>������̧ť��W>���oq� �w�W.i!DD*��!׶.H���z�2�4��]�����D�Y��.F�<��i�W�?�?����@

��̀�'$Vj�����q��J�U,��4pX�JOls�9 �]k���^ y8������K&'�^g{j��7]7�\2��}�S�Dy�t��_M�M��jG�d�t����Ʀ�0��Z�zkf	�J���ڬ�ѓ�o/�n�Lq���8s�5����Iɒ|[��j܅B��5��0��e���	�ő�d�4�Z��o����8'����;��e��r�ҹmVK������yKD�-#3�,�O�R͆d����D��|5'����
���\����HE�΋E��~GJ}�j��O~�{�K��!��K_��:w�/ll?���(��y��*�Si���K��	�b�OPюQ4*�F`p����ƞr���x�w�l�EO
{��$���e�ĶsG��t�ˋ���#�Vc�B��h�N�"��g���|c(�:Ҡb�c�Cf������F����H��� D��
�9s�G��z��o>h&�U�9�_��c�$2�����]˷)�F� ��R�0��^D�	������K�i%Ө��LR.dI �:�Ǚ�oג�<8�ؔh�|��mP�䟭H��T�/��NH�vI�����8̳�Y�=�I�\K�L6�0 �\�Ʋ�Ɔ���W�M}zMW�x��]�6�@�m{L�|�٥��2�m3�Hw0�6��{%���Yye51WZ9v�Xs�q�����*��V���.0-ϴ"�L��9�y��wU���#��[R9�]�R� v��zB`�����7u�p�M�K�8� ��;��!�2��-)CX6�E��$��W���}Ay��{> �Q��yC;vZ��>�SJb�7����m��n�N�l�)�x=Ky��O��1�L�]�Ԡ��n]�k)�!.h��>��i��ꎷǔ	�;c� �b~�~�2$�#nptm�����]�8Tt�&�Oo;�����.غ�5��5ÎR9%�g�O=Sk��O��b�v
�W|�4kL�"��1'����Xy�uS;�/7�=����M�In9���uM'� >��'�m<% ����f.+I9��jfG�[ti���д�v;��W���,����d��n�t�Ʋ�F��;��(�e�MK|g��WT�E��Wc
;&����6MGt��s�Q�5����*C
�
l�.�L	y�w��"��2���h�~|&���2%���xp��A�F`�{��f�<�9/��^SA\������*�R�L�a�����Qi�J9��L+s'�E}	v1=*Ik��Sr%�	��5��^$��E��h�8c����%�����޻L~�HD�}��*YhW�NI��b)�Y`ݺTd!��?n���s=r�q�h;(7YC�9�m�pЎ�.��dhW/M��iO�o���_ PK���0  �	  PK  ў,J               233.vecчo��߽U�D��*1Klb�FbKԎMlb�c���޻6Ե�y��䓻��r��H
#q�(���ԤEԶ��u�G}АF4�	�4��iAKZњ6���)��䢳v�+��N)=�I�$��ڇ���?� �ѡc8#�(F3&���:��1��Lb2S��4�3����f�ʙ��1O糀��/��YKt)�l��
V��լ�
c��c}>���Mlf[m��vv��]�f{�g�_+8�Aq�#��q=��$�Sz�3���,.�E.q�+\�׹asSoq�;��g��<�y��y�S����^�����[��|����+s�����o��=���O~T�o���,�PK8��c  �  PK  ў,J               234.p��y<����c�a��hl5c=�%c=cˉ�s�9a$K":Ӑ*Kd?v:�$�d�=�D��}92g���?�r�}������|_��y?���aOG͍͌ @���#�������7�����OLP�J�8��q4ZBF	+!� �F�N�*(����a�ZM����~?�@������%ђ���؏$7H�I`$��� ��'�Հ��¸��^΅�G0C!0��s� 	�T1�"�¥�(|ԭ\ni��va��2�n���c"�b�O���d���5Nkj}g�=�������������ٝ�q��wХ��ˡaW���Ү��ӓSRo��gܹ�� �����������o��MO:�O;�XϺ_����ѱ7�3og߽��������������� ��ۿ�Br��P(
���/�_@Ba�*\�$�+UH
ō2��[ݎ�V��,�8�sLF����}��d�X��D��r�|�y$�|.��]�9Dj�#��7b�ڡcu|�Z�2U���}{�����V+����@��MIDp�@�T�[����
 �E>y��Q�󳉆p���\��duEA/2��\pj��Yl!�J�5%ƭM��.���^\� �����+���T,��.�S"hg���l+U�c��$"�
�o��V	�Rfьd��I��2����O�~"��}<y�d��h��!*3۩--��ͽO��������w�ľ�z�q�Q���7�Ȏ��.s
�'D���9ԑ���4J�[ %��,�cOR��1=�]�I�5=�T�L�	�un� ��yb�8�s�7.��� ��`��	*
�L��Ud��U摗��������θ�6%m��G�eQ�����C��Xm�_ȣWǢH��$���X�$VNq`��U��]ϯkV1���mW��k�S�ԟ���$������/.��M�� ��̚	Y��
w�[�Q7N=I*EE�4�>��_���@s��+��O�m����͖Q:�\�6� ��Lw}��O���ZP@&�Ӗ�RК*�O^�{ټj��u�A��c������Ew�w�%{��V�)Z�ؽB��Y~+�,q�a�VᲮ��4	�)�E�Rj��h�_"�g�ń�ݲV��ɳ?\�Q����5�����e4B:*g~
�L[q �u�m7���G����:�70qJ$[�ai�X�R�&&��gؚ�#�����ū,�x��6П����e�\�cO��_�y^s�F�؀9kF�Rh������i�ؼ�������k�s��rh�CjѿޯU�����g��Q��>���	��7Y�S.��� l5j�i Xm��1����A+�uZ��%E	g��V����6��E�)���sc��&����*���J�]��l�O/�Cc8*w(�|f=K�Dt���_�#Ž>h5a�
L��j�[��#!ɳ7��=��צ�/��f�P��*��k͹��S��R�0<�Da���>t,E	"$�.��4���k߂K_����\�8���H��rbBQ7e�=�q��D�@��`\}k<)��jV����xZ�i"�.��� ]���eD�j?~6��w��̍�
a�Il��������8VO�eCr(e�u�酽
�M��N!ɽ�B��_0��~�<t\)����Aj�eM�Y)���x?�Ȁ _1y$r�,��h�^޲�X� ���b�?*��쫆FΝj��\;���%qDƗZ3tjã����	�ˣ�2{��3	��O�l%�DJ{�#6��:��{��م�*����a�v6�n�3Q����;,�bw�y��In����{fb�VZ�]�ꙇ#:�@��&�cph��]vI�������o�G�PKF7�h  '
  PK  ў,J               234.vec���Q����k��$VM,��Kt��(�D��jt���D':щ���폚u�#'O>�ɛ�ˉH�"qr���?5�E1�m�h]�Q�4��iB	MiFsZВV���6��e���\t��t�+�(�;=�$�K{Ӈ���?� ��:��c8#�(F3������L`"����2���`&��Me����<泀�Y.�b��,�e,g+Y��j]��B�t=��&6�lѭlc;;��.v��f��c?8�!s��6��8'"��z�Ӝ�,�,��.r��\�*׸nsCor����;��}�<�G<�	Oy�s^��7^y�׾��w����S��Ϲ,���{�E����|u������PK�^�V[  �  PK  ў,J               235.i��g8����,VoA���H�w����A�V�V�aW�^�K6:I���`uA�²���\��9/�9������=s��\�\-�zZ�Z 1 ]�jP����d��`0��������������;������G� �~NN!�;��$%%!�rJ��w%$���	55+�8/'���s\��D�\@�@b �� ��$%�� �G�HH����T�j�b"��DJJBr=|=�0�2򊩒�0��y3��%��ۘMG�
H���)(Yn���ߺ-($�������W�������3��[X>zl����������+_?��ׁo#��c��&%�������_PX������[uMm]}CcS{GgWwOo_�����������*fm}csk{���{���w�." D�?����p�ELB"������?HHy��UM�v�7���ș���m����ᣔ,�+�����d�w`��_d��s�� ���1 *�a�9<s ׆�&�&R�M nO �����@S�?/]�z�5�CS��~[�v{>�hH%�;A��0sۿ���4F	n��V�l����|��s��|"O��$'7����j�*^��J�b\Q/8��>\��xQ8��xR�Jw�rg��c��K�`y%X�$ډ��ח#��X����$1��a�!���hZ��!i�ޒ+Xp�
8i�a�]�tAP��$�4F.�n�d����h���=elR8
�M�yg?%�Kt��2�{���2��vؐڻf;GLlV�z�ӃÖ	�	����^x��\��V���P"�T:�~�'�apS��_`3������f�(PR_�)C0$�ip-��iR���~qvbf����2��oyTdOw(G(�Vb�D'��V>�4��@4��	�фHT{���>�*���Z����bH�oUu�	�1�Wk#��at�\�%������� ^��w��<�~̃���R�x�:)	3x�A�A-1�TV��5�sJ�c˴�uB�&9��1�7���!�{�ҋ�֗�C5�<ymO&OӉ��OV�����Vr�h�?�?I㨎��rW��Qq��:�yK_�U.>2���"���F8U�
��aѢ%�s���p~����&�
��.����C�Ԇ���<�
��i��Z��k8ǖ��Hw󞶣_��A�Ez�۝�{��s�%�u��d=�'���4��n���[d�i�y�	�L]������p���G]ȝ4ђ����`w��A*��W��h��IeY������~<?}�ǅ���s-vʡd���މT�ʻ���a�f�]�a8�u)�˗Jښ����l�7ydijj9 �</���ĮyG�t�����6�}�R�($�)�V$>1ߝ��,�!7�n�����ex¬�L�����j�����F|���w@�����K�-�&+�|,�ƈ�[Y��e��]��<��S�9QS5����:��o���,��48y& dC�Ɏ� ����܋eG�M��3��1ߧ�bDw���"��*�
�d�@�zH8sJHЗ�#���Bw�2�*�Y����v��T<=�S��SfL�o<��V9CP�?��m2nF&�u�T?��y���
�*�sjp1:��~]�e;����B8�Tԡ"��c����ɾGm�`�OW@�<�Fs��Zԃ��I_E�i'����oⲹ�
L#@��y�����3��.U��8�+���i�����4=~�c������N��iv��`8�L�m��d'�߇Lb��z�V���D)(|MIqFٵbe/�"_��m��]�J��#��WA�/�sBj{=�o�!&?�� (]'5Bom?j��[�+��v<2��K=۟3�>EF$wPڱ~�7�í��lK���51�����E�E���
�z�^��RI�'��iR	��.����d��f�Z\1��ب�X%�g��A�p:�|v%Y�p�m�g[-�v˦8����{���ڧ�Y���
gAC���U*ڽ���'x��h_�n�0V���1!�y$$���$�Ơ��Q�%_>/̃q�Ml�m+z�D2 �8����JQ�d�����+@�cH!���Jx�2c������\
>+GvV[�"����1ߋ��Xf�#�ʼ���	X��+y���m[��y#ӓ(���`�e޶��㰭�PU;/W�%� ����Q��݆���'r������M��q�(�Ǵ�BR�u݆K��ؓ�o�73�5c%��^���݊2Zuӈ+�WP�_ҽ���*�|�<z�s�V1�%���}��X2��z�����	d����@ם�@�:(��3��o�.��
>*�8u,�#�"(M���HQ9��y�h�:�ɣ��y��ɇO��8���K��C?�9P�?ߧ޻I�!R��ʉ��a�-E�b�yr[BthC�:ȔN/��c#s@i)�6�G��)s����S��Gp���1i̦��Zb/��F-E����~�e+r#҅��H9�'>��(ˬ4�5�������K�:�7�����@�CR��r�K��~pעb[�P���Ѐ*��p� 	F��oC��-h����y3��ɠ�G]��<o�+��_��JG��q��{�[��N�G���x&�B�nm\rX8��`"/[IXEGm�h�����y�}��?+�;n�Q�
_n�>���u�4?��Z/a�]^�-�w3�_��T�d)n�E<��tT�� 9z�o��;u!"�ڲ��ٙ�1����U��[�u�wo'8��@����Z?�!�r�UWx�ᾢy��!�W��P9㖩g��y�=�Y*���WMFD��?j�Fn�[��դ���-ͼc�ˁ4�)�� �;�&��H�Q(��N�y�	�|���!+`,b�ri`�����/�x�=�'�us�X
�������t�_�TƎO�pһP�����ޏ/�]
?SR��R[��n�\��Q��n��đį��y8T_S��N��]��c��fN�y�������[##Au�M����xvT����N/Vg���(K,��Y��$�����e�}MW���K��S���H��<���Ҋm�W!��Г2�`�k�+�75�y��s܃C��]���h�Īo]�[��O��8�nǵ'jt��h)�Z�
M��>�4u�%�T:T�q���{�����°�z��K1X������(��Ή�,^�"D�@5ƶ�pzT��_V��l�W�9�s%�X��*��L�c� I_\���7�*'Xk��b/��/�����݊�[��ǺNɊ9b�[~?U=)I7��m�x�Ю�/!9a�A�Z�#}Nmw^����ZHl��Q\m��{�&{S4:���n刯 ����ަ�Or�L���[�C�]�6����i��m늃���PR橀�}��.�ٙ�Y�J�i��N��o�(4���� �}|q�w�&?y��v���ܺ��2g��UAy^z�总���l�|����� �?�'�Dփ��}��JP�&���V�a�@�5(S�����r�.�g��� �$���k���]17��S��a⦂�]W��=�L�Ɗs0Wx�!�q�c�m2�X���"����.?�1޳�nX�w�l�}F(��t�kNq�����I�<Z�~H�ъ���M��FK����{�F����Msh���jN�SV���F������$�Fc�S�cp,[լ��2A�1xj�,�T��:�@�@�-j�Glmy^��*�� �����U���YiLy<����z��6�y66�a�����6j($|n��ž�7zs�T3����L/ЋLEoc�*�k~�t�۝�?���3�L��A�5ki%�de<��9�:��y��jС�zv������/n���D�#�<~�f�sm3�-�h͍�DԮ�d+{a�2��nHw�|��V����j宀��}�/2ن몠Ep���tZ�0di�n�\�V-�cq��N�BPڹ���kK�I�)/~���p���aύ��`w����d*ektVi��|Tq�����Xf��̓:o��:�N��BL�����aY��oz�����^�d���/��y�A�	D��-�[b�,�/�Z�
�H>����rd�ۣ�X�O���r�Pf��wa;�.�U�=9s�5=�y�m<��A�ԅ��k���<[��"~�[�5gY�{r�����a���z�y����RңM��î+��Rs���|�h�����+`�J4ąc��x�%�	�|@�vκemC��V�����I�LZ�ۢ�/�~zt�D�S��iO�����,�b�۽��U%���~%.Z��|{u�[�}5�d��IRN��کiMZ�`�A5�!zNv{����*���q.;�%W �K���2v�p�H:��[X/��M�"aL� �Nݵ���k�獛*�~a{wC������1$·&��԰��5R��� �h�n�����$��~�^�X����	��n��9����q-���򦄎�@,�h��v�����i��z�a
�1
y��{ۮZ����̒%Sϭy��vS<�c��G��{W@vj{�a3=Эo�mu���/nqV���ij��xtW�fi��Q9���)L�O�i���{?�~C����r��r��v�tx����@T:ŗi�ƢG��S2��0�tR&��WL� �{�ۥ���6�}��ʌ8��4I���e�U1̙JZp�/�M�]i.��/>��`m��oMf�E,�a�xm�l:�޻��P��C,6�z��R��g���0��##\ˆۙ�Pф�q�����|������ÎnYA�^�ݞ�&
nTEե�i}>�~F��\�,�6p�
	fޚ��(�5��u��]n@#��V������a%i�t5���낔k�B������g�@�)�;��?��~�}	��WJ*ʻkd~�V�zL���R!BJJ��1�4%�F�Y�J)d,�s�R���լZ.�S;���,�n�v�8��2�O���!���<���-3_��]K��zc���j~���e��?Ր�������O�T�2��®��["G�p����";��p�&��8]M�=��>�;���c��EmuS֬.�ด�nӈ�C(������-�Ĥp�:�M3���)G}��<�����6�"�H��cKf����>�\5l�p�
�)�	k1@j�����,��ZE��N����������Y�,�{��},W2�o|fb8�٤9"<���O|O���ҧ\3����E7���d��>D[�f>��i����O�C)�W�����6�x�&�Ues�$"bX/��}�}
�_x(��!я���m�g
�|��Y�_o|c��?t�Д $-W0��Az�p��|���[8�9a;>�#�*Ûƺ�!W��#��w�y�:,�]�R ��*η��s�֮î��5U�t^��y��G.Cr�ڌ5z�y���N�-��2:�0�%O)�*�Mkє�9J���
�vW@���6�Q�w�__6D�5���gu���+#qW ��%<d,�+�����ZkY�ځ�5$%"�F-j`���燊s�5-��g��CյL��<+A��t�.�E"#�rYff�,[I��:Q5���P�R9��u.�N�Fym�e	|}��z^���.��~"�P���L��	�����Y�ӳA�e+��4c�w}Q�3+�U��u�8G�p���ᰕн��A=1��l)�ߋ�0BjZ�o�"���z��T(�β�~��2.y����y�3��G���&c�(F�$v��x�L�$��"ϳR����)b���\?M�˓*7M�"���(��*��ԔmJ����Q��лJ�Y�������B�G'��O%�r�ٲ�����>��I���B���ɱmP,$pcK8W���?_�>$��*��A�)���b��'�s.�Gy��Ja�2�b'��r�HY%C�� �r��r�z��J�x(g1�o��W�e�I��a,X���2��$�g�=8|��[S
V��ӏM�?�?ɫ3b� U#��]��c��7���H��ｧlir��zI`sR�!���}d���������]�2�]�v��Q㬖O�ER��<��#)�m;"bQ4���Jcѽ�%[>�'U~�mR��#�B�B���p��	�\*x��$C�;�xf��C��ǭ����+�/oƺU͒y/ת�H���:�
S�9}o|�%���l~��*f2Bd�f���U�&�{�KKe�ȼ���q�Z�؝�Å�C������;>_
1��h+i�>,N�!n����Fqi3R/�F�EM:��=��,s���|Ӵ2z��g��v�.�Y_�4�${a�|d*�jǯi=/I܂��9:}�>Ǘ�e�W�2/�9\Ф�,|�!M���_�Y���1޴k��0���4�N�@�����۶���삁��/<[���|��0X�xVP~羸��Qx��4��%�����fJU7��/9��L��z��\F�!q�RIߔ0������h�6�+`�$~�iJ�_xm����Pq��l��9��|r�3�pz�F�TI��b4�E�����X*��=f�;����O ��^�_��ʴ��$��<�K��d街�ǐgD�s�[��ے�n�q��j�S�9�.��x��1���̿d,/�!W w������ܼ.�ec[kU�aˣ�qԝR�ʡ5^tN�^����I�˽�'hj��o��ܾ���.TC�,�q��R=����ۻl�J��������5ԙ���A�d�0��q��/%ZM�uM㯥��������g9��W'�L<����F~�$��`s�<��d������X������8s�㱜{�����ג�{1q��gW@N{6F�=�k�	������2]���]
��O��uĦ94�)`�JRB���J����.fڸ�
ci�]��U{+Y_�2A�Q����8"Z����a��Yoe�1z�^r��=�#���`N^[c�%=��@ː*8ݶF�Ob:s9B�X�������}�V�`���Z�w�r�珋FS�]H]����ܷ��/}�*��q|�'l���B��;���tf��>{h��^�Q&N�Δ�kd�k�N�[�r���F�3�(C�c���T��,�%��3z�-iRW����!�a��mm�Q�wxR
���o���\{�g͘5u��7H�|�����c'�KY��?��0����kQ�9��-�Bݗ|ܽ,����nŜ��/��DHV�T#2�
��te&����=)�}&?��d�Ed*�#6�p"ť�y�#1YMTV�h��(�hǵk`Vg/B��ʼՙ�G��L|_�!��=1���FDw�b�
��ߨځ���F�mCʾ�W�M��jL=g���ka^�J�ۖ�u���<��܍��N�I��6�[/�v�;�A�#�u��cɒb9W��PK��A��  �  PK  ў,J               236.p��y<����Y��h�p,�h��؍�D"�#��e_�(I�(e�6ٲ��,��F'G�h���:�T�0w��]����}���y��z���z����>��7�[k�5 B  @8X�bb1�8�@"�Qh�$ZB-/���))(�����o%�l�J�R�����Zz�m&;���P��7�H$Z-'))�O����6qpP� B1��P��Q�?
�@ap1�8%!Zpw �P
��`��(�< ���	K1,�A���\)W�ͽ/�c�<��{:���^N^AUmY]����x����_h�{l趎:9���>���X���0f����q����Y�Y�9W���5�]�Sٍ���+j��r��������������������C/Gߎ��'&�MM/,~X�����˺@���� 0�X�!g�``pELڒ��	��c�q���p�#U�?�����EɒFU���0�6�����_b��z	�������� ��Q�`t~����v$ }_(�y�X�
���7�eH�����6�l �|p����Չ:E^�����(k��e�L��f:�A���k���-/Q/�C��W�V��y�����y���p�Hi�ٹPt�	%����q�_<���,��ѓ*g�8�9�d6��c��	JU�Aĸ�%�;|V�!�E4��5*�aA���8&Yǋ.G�����pu�qm=�3�1� ��˳�s��ȶ>����5-!@� ،��޳�ei�h@���!2/v�P&�4T�����Fo����n�$����z������t�á�_q���C�����>v��J�Ƴ4����յ�eם���=�E�M�%����t�˩kkl�Fx�+�<�һ������nD��ˢ���4`#��
̑|{)9�t@a��(;��L�r� �do�����B�Ԕ�mf�RRڤU�l�Pm&��+ZGA�r
[�?�a��8ѱ&��������Y��	s��,�B��M�j��^T�����ۦY���#{"��yYN���h�i{�=2ol �ERaz����*�'oC���X�:�`P���d{�U���M��_������.�A}�QG�v^��7�	�1/=��K���Y��Q��W��55k{��x=YM������Ot�I)�/Қji����y#4��~�d8�ǡ���Q��`@y���T�aMk1!0�,W� bZ�|�ǰ������p�YYj[_暤��punU��U��=?�xK�?%�,�������A��/¤�*ʽ}�f-�4�o���7C���YO��Z�\ef��a�\�]�"��˂u��wv�|�����o�+�1�I�AXb��7�Ԯ��g��.�K���X�c�j�=��^�y�x�E
WW�=y"\�5:e��ġ:�����5}�_M��"W�E�����i�?�����w �N�Ks���ۺ�r�-�rk9����av�#i��}���|44�<��ÚF�ʤ��C�'�${�c�clVM�&���Ҍ��ӕ��i��pD�xڼX����t���ecU�x��H�\���=�t˽�C�B h�~f^C��b+��j�t|h�e���yJ��Է������'�#�%�Q�*��G��*����;������D�Y���������t䍲��LPVgmR��c�m��50�!���f�c��^g����T�@uf���`
.]I�~{Rt�S+8��d
�� o��>7��u�u�#�ډyW��v!я�"h���]�na���w�Z2�آ��h��F�S��yU7j���¡�PKQWu;  �	  PK  ў,J               236.vec��ˍa���}�ٔ-�l�ɦle+�l��&�l��&{���s�sy�����������E�ˑ���T���bSU�Q�Ԥ��C]�Q�4��iB�,ʹ9-hI+Zӆ���r�^;БNt�]�F�,�ړ^��}�Gd�����2��`$���2��L`"������S��tf0�Y�.b��e�Y��E��%6Ku�Y�JV��X�kX�:ֳ��lb����6������j�u��^��~p�C�Gm��qND!N�)Ns���K)��.".�e�p�k\���7��m�pם��>l�#�<�9/xY^�W������|�#���"��J����=��G��ɯ|1~����?PK7��`  �  PK  ў,J               237.p��y<����Ϙ�C�fl�Ӥᘅl�`�dr.�B]�5�,Qr1���DS�AG%ʖ�!Ke�Dt�Π�f��u�����������y^��y���H{������.;  �l �~�@��8�@ P(�'�A�1xeEq��q#���k�EK�B"�۷R�Cs�����A[��B�0h����:M��M��KZ`� +�*��� $m 4e焁����!P�Dɡe*� 0C!0*�=%��X��6�	W��!t��h	Yא$�zU��]�X"JNm�:~��o����1�������ز��v9���s����<x����Q�1'�$%�=�r>�B�9/]����F���[��{?WܯUU?~�����򴵳����W=�}Co�G������جxn~��ťϫ^  �G�[/���B��U/8ju
Ӧ���qZg�u��E��̨��uȩ�2�6Ϯ�}5����'���˫�@@�˃`K`F@��˭���.��K��#�d\���+�܏����
>Tp]��ʐΑO=�4�޳�$��Ѯ���b�>�o��B)��neJ�ԅ�U`�����2ΕL��XE�ru#V�>��E��	��a�Q�E���oJ\tj����b�>o���٤����������r��=�JȺ�6��kj����5<���[�?��Q3(�3%��>F������&�.e�qwC~*� U���o�٦�B�n�@��<� �n�T�ӈ��̶�z��B�NG~~ڃ*�>�����B�w�o��n�wTg&�xy���C����sa`1cj�io�H��&fmO\�P�&W�69�����p���ſ�Q��$uuWZ��T�f'�E��Ԕ�^�l��У���|	>�L�d�*��>��w����0�F�ٚ�YiA�v��܎�8�"=T�WM3�[���)�H�n-}��)I��d~I�z;���=���6(��F� 	w�QF
Zꍮ�gT�hSW�}d#F}�v4��.������9) �Z�6�����ŕܱ�e��Xs)#<sxGt܌0��b�z2(�۟v֋�1f�bĬٌ�u�]%5Β]ES���v�L�/��\�υ-�R�No,��e}��Έ����w{!�q߶����F�թշ�x*������ﬃO�	���þ��馟;��Cd٬�:$�ѥy�(��}�$jG��U%����'���=9݇�SU�������[.;�ѷ6y��5%\���-gu�ŜG,H��y�\��g��fw�pM8X�H�ސ	��I�ҕ���w5���Ӥ�:� ����R�3��'[��?����[��Sdos^﩯2]Q$�W�s�tpzGs�	���j���}zV�e��m����X'�.!TI@��7z�.{E�q9��������c�ؠ5@\���^)������c�z;$�m��?l+%B���Y(��^����~��c+t����>�T�:��xRE1�X�,�u��H|lPXD��/�!nr�\�<-ЩNK��SP�og�xɮz�5+��U�2u�U
4�Z�.>�C�uE4�R�����񍶵:~/9�����S���/7|������M�{W�e�3���Ҁ�rg�id���(�Zs�4��)�AS�:�����&�uϐ�nF�O3&?�S����^h.3ü'�KOΔ��B� _y��͛�@`�R�w�J��`�0j��o5��J��"B�Q�z����\�r�����1�#α��0�EM�q�`k��,O
������W�B6�sh�d�f��6�3�zE�i���B$킩{�`���<��Gw��^�@�2S��QJv��.�1�P\�k�EkA.�6N�q�[�M�;s���md]X/��7���? PKU7�q  ,
  PK  ў,J               237.vec���Mq����_��*[6�d�M��V6�d�M6�d��E��{�Q׽�=O���pND��̕��J�R�*T��)�5�Em�P�zԧiDc��4+�fڜ���iC[�eY��t���BW��ݦ�����C_�џY1� 3��c8#�(F3���c<��$&���S��t_i��d����s��|���E��%6Ku�Y�JV�|��5�e���F6��f�ne���Nv��=6{u�9�Aq�#�9��9���I=�i�p�s���).�e�p�k\O)n�Mnq�;T�B��{ܷy�y�c��g<�E�/��W�_󆷼�=�ȧ�9W�/���չ�R1�G��̕���O1�PK@T�9c  �  PK  ў,J               238.pŔy8����/Y,!b��ZB����	3�j˘��u����f(��R�.�K�Ҫ]���֒Z�j�D����D���s�{�y�����9�����9�7����a{  �`�!�B��)���D0h4FVBR'/GP����U�5�����D���t�&�$sm}��!$�AcdDDdHJx%���f +�n�e ���X� �C��π@A\!�D�	U� �P��`��3�} ��K(��IRʑ8Rrv���my��[ϼ�~ =���##+���Aܫip������� ����aG���^�>�A�!�B��8�CtLl\��s����v�"��̿��^�c�����݇�U�5�u���������[狗�}��W�co�'&��Msy�K�+�?��osA ���\Xa�m.4v;�+�	I�P��ʤda�mv~yRE�m^*�ރ�V5S[�F�B�����)����k��A�@,`��%��P����`�g���O
�Su���'S��(����I���%�#���~��T�T �S��O����ke^��6ɳ�FF�+�I��Y�lȸ#�?� �d?��Ac"�&.�J��ng�0�sS��'�m�mՁc��q��l�M5g�	I]5� ɎvjP$�d���OM,;%�N�p_R�>��ri0=�-�`��9y�M�@^d �@�y$Q�8��˛C�PU��jki.>[AKl�_>�	{�@�8ݱ;;��9��3��T�l=MdU,q'���'���{�`ծ��5/����e��j{Fu�TO�].�G(nձ廃`9��<�Tf�Z����S�Q��B�����T��갴�51y�����kT��I{B	)$5����$r�J�٩_Z��V�]F溝�M߉&����մ�>�=�knwF���>ɚ���Ԕ�u5�Df�j�hK��W^��8*�I�7���ǅ2����A��a����KXɂ��d�+ħW���r�}�L�1C�;�}_����x�z�EpmG/��=�Y�S+�e:���)�[Hh� ڝ{)r�K�.�L$��~4�j�δ輮�bh��T�����hc�e���y*-���Z=s��G,����ˍJ�8�9Ɉ��ʆ�-*�v׶��Y��c{?�8�Q~���ʙx����(��<�Tc���c���t�QJn�d����L�6X����
p%��m���J� E�&��
Ĭ�ʧ�5�3S�w��9f�*��������f�@��+[�v��~B1ܨ�Guء簼���7Reo�f�yv�4�A�dλϦ����l��)�+���@�ZEΌ���y��F��Bb���-q<�f����
A��X�URɤ�6t���o��;�%\j�B�V����1��a�bK&WT-�{��9�N���"�������@���C���=d���~6�E��`�u~����]හ�=�ok�P�����e��d,P�s�i���ݬq��+&�~�"ߛ��phy:�}�b��#1v��tStl����k�VA��g�ee��'&m��s��6;�+��1>T�=\@�Y�Ӥ���"h�/ny���!�:��D��nE�>U�Bn���`���6R'�G�_)	�Xl�K��&�뱯��,߷~9#�5:�5Q��&*ݥ#
�1�$�	sӚ]?r�`�l�NPNO�'U��8���;�b�mA�s4Gm�'|�N� IK��M/�f�;+1��MF~.ߐr}G3\TC�����9�2z�,-��f�8K$�U�P��y�^*��u��v����/7�QU��3���w�k��j�����5�@�A�U�K%�g�)ǵx����ѿJ���PK\�J  
  PK  ў,J               238.vec��Q��3�]$����E':�It�.�%:щNt��(���w?j̎G&Oޛ�����Iq$��(����Ԡ&��M	u�K=�Ӏ�4�1MhJ3�SJYR�ڒV��miG{:x��ډ�t�+��Nz&I�����/��� 2(�b�a(��F2�ьa,��&2��Laj��4��f�K�t6s���1O糀�,b1KX��2]�
V���yq�ѵ�c=��&6���V��vv��]�f{��������9�Q��9�'8�'qJOs����|���ȥ4��z��yQ\���0sSoq�9��r*�4��=�y�Z?���<�)�x΋�,^���k��w���d��I_����<���~����O��PK�2̺f  �  PK  ў,J               239.pŕy<�[���1�\#�\[k��r���2d}�l�0e_�I��yQ��U�ɠ�h�VWȐl%[$f�t-1E#sG�g�����������y�s��������8���  0 ����a08LH�#�"��()�O\B#/�𭼌���~]uEem99����A�@PP74%�Mt���E@B)*�BI����u�[ �0��)`4����9�@_�G���.�A
&��� �	A��l� @�B�J8K�����'g
�X1K�,���LA�앒�'������$�2 }gM����wp=������t��	jpHTtLl\|��ԟ���g\��\�r5���k�E�%�ݭ�yP[W�������I������/��GFǦ�ٜ�ٹ���V>��q?~Z���� ���B��P(
����'��BJ8��%�!��O�Xe2#T�\�%"D��'L��l�}%�k`)�ٿ���5�B@� h�X��e��EMVɕj�%R~~��q���m/�0\��P� ���=և4~�T3ַ���!,l�7�>�2�N�m�%~?ƞ���y�e{�GbV$�� :��3���D�aZ���&!@�����(��tÆ���x!�D���z֢���rF�Wxf�Ew�BDO���MQ'P����^�މ�!��'U�ߎ��q�|��y���V[��#�?n�Y�Sc�t�?h�S���r�A��� 5+���!X��������gIUoi�a͓�K��1�"ʬ��f��Ds�
�<
��iē�52�
"a�w<j�Fe^=SB�R+��aR��6�����!��$�g���"J��%���Ř�E�O��*eЙi����O�Wݹ>/3��;Ǫ��xv7��,mRh���:E�������\�$rJMv<Cv�ɚ���XO"�? e�y`l�G��<�ý��ҊW��+f�3�S׀��()�ƫ�ʠu.0w��f��)�|+{����g�~���+yB:����L����%���f�_u�A�Id۟��3�At��H�Y�uw��%.q�#0n)f,���N��v��^Kl+I�]s�w�	�1R����E�u�o�e���d�%9Rsa6�����%�Ir�s���^D�N����Z7��)�ߦ�����yE�j�C=4�!f�ֻX�z�x8��ɚ󙸜�v�<z��Hp��ܽ�\'����� I����2f�M�Pf��+�{ɵ.w�Y�>s������I�gtE���D9��ũQ���7��v\�a���A�,�E����N��|�(YԢ	�*��飴4��s�����WĀ����1m|��x˓ӰF�k�j&��Ѽ�����phR1�ЃE7�`ȇ���]_;�?���K��AW۱*ݒ(�S��|@�3"������_
:Ӄ�tmg?U�5�T �;a���l�%u�s7��^�W��c�/Z|�'6��R�p�S�K�Y+A<�c��z��:�X,3�@b=�R�B�
����t^^j��ۦ��zu�n5\c���>oѢ������e�Y��������A�ى\��kΪ�ےIRk34�w�̯msK�|�Q�3�P=�+��3GB���/���H|S��+ۢ�%��O�07^�c�,�:�gi�C*�������2�@�F���Ȧ���������
����ذ��|��x�J��:�c�@᧳J�lW�̼�޽t�],�Av�W�w����:���V�\�\@���Q[�s�6��.��ț#�G?8F��d�gUo���̆�Lyd�x�X����w{#D6ߘ%���QaIa�ܧ�A1�&g�J�~�R(�ZV�+����(l�P��3Iܻ��=�Z�������9�PK���C  

  PK  ў,J               239.vec������}|�([ٲ�&�l��U���&�l��&�����Q�>����{u?�]DR��@���R�JT�
U�FujP�ZԦu�G}АF4�I�DSmFsZВV��m�b���t�#��L���s�kzҋ���/�蟔b�d��P�1����Q�fc��q:�	LL������T���tf03Mc��fs����,�B�,�%,e�Ya�RW��5�e���F�M��-le���Nv���=�M�ا�9�Aq���X��q=�INq�3yg��ӿqA/r)/�e��U�kz����Y�ѻܳ��z��!�x����(e���|��5ox�;��|���������g˳����#��Y(�/�͟,�PKt�m�h  �  PK   ў,J[���2   3                    metadata.datPK   ў,JM��"  �"               l   0.iPK   ў,J	r��  S               �"  1.pPK   ў,J,�5�p  �               �'  1.vecPK   ў,J')  H               �)  2.pPK   ў,J(�l  �               �.  2.vecPK   ў,J��{  :               0  3.pPK   ў,J�e$�l  �               �5  3.vecPK   ў,J�|�C�  4               W7  4.pPK   ў,J�)V�n  �               �<  4.vecPK   ў,Jrj��"  �"               &>  5.iPK   ў,J9➇�  ,               f`  6.pPK   ў,JI�x�m  �               �e  6.vecPK   ў,J�$j��  �               ,g  7.pPK   ў,J�Xx�r  �               l  7.vecPK   ў,J���  �               �m  8.pPK   ў,J� qp  �               �r  8.vecPK   ў,J��ܥ  �               3t  9.pPK   ў,J�Vpp  �               	y  9.vecPK   ў,JS�q�!  �"               �z  10.iPK   ў,J�g���  �               ՜  11.pPK   ў,J�{ݘo  �               ��  11.vecPK   ў,J���Ԩ  �               Y�  12.pPK   ў,J�o��q  �               3�  12.vecPK   ў,J�����                  ة  13.pPK   ў,Jl�&p  �               Ϯ  13.vecPK   ў,JI$ٸ�  �               s�  14.pPK   ў,J�{Q�r  �               J�  14.vecPK   ў,J��B�"  �"               �  15.iPK   ў,J��R�  �               A�  16.pPK   ў,J���s  �               ��  16.vecPK   ў,J�� �U  �               ��  17.pPK   ў,J�@�cr  �               "�  17.vecPK   ў,J��B  �               ��  18.pPK   ў,J���p  �               <�  18.vecPK   ў,J��]��  _               ��  19.pPK   ў,J�M5�v                  �  19.vecPK   ў,J|6M"  �"               ��  20.iPK   ў,J��ɕ�  I               � 21.pPK   ў,J1�y                   21.vecPK   ў,J!�Q�  P               � 22.pPK   ў,J9��|z                  � 22.vecPK   ў,J�g-
�  Z               � 23.pPK   ў,J�#_ y                  �# 23.vecPK   ў,J����  I               |% 24.pPK   ў,J��w�v                  �) 24.vecPK   ў,J �p�#"  �"               @+ 25.iPK   ў,J{I���  R               �M 26.pPK   ў,J��+Pu                  �Q 26.vecPK   ў,J��K��  S               gS 27.pPK   ў,J�@��v                  �W 27.vecPK   ў,J�d�2  �               5Y 28.pPK   ў,J�h?�w  �               �] 28.vecPK   ў,Jٓvv�  P               D_ 29.pPK   ў,J*:��v                  dc 29.vecPK   ў,J�I���!  �"               e 30.iPK   ў,J}��  q               ;� 31.pPK   ў,JI�0�y  �               r� 31.vecPK   ў,J�_6j  �               � 32.pPK   ў,JF�i_m  �               �� 32.vecPK   ў,Ju��>  �               \� 33.pPK   ў,J�귁o  �               ̗ 33.vecPK   ў,JvuTY�  �               o� 34.pPK   ў,J�(��o  �               %� 34.vecPK   ў,J�3\�l"  �"               ȟ 35.iPK   ў,J�.
�  �               f� 36.pPK   ў,J����l  �               � 36.vecPK   ў,JY:�_  �               �� 37.pPK   ў,Ju���p  �               K� 37.vecPK   ў,J_K��b  �               �� 38.pPK   ў,J�$p  �               �� 38.vecPK   ў,J��?^  �               '� 39.pPK   ў,J�fU�n  �               �� 39.vecPK   ў,J�(���"  4#               Y� 40.iPK   ў,J�T�t�  3               0� 41.pPK   ў,J/�&s                  1 41.vecPK   ў,J"�{�  M               � 42.pPK   ў,J0o�r  �                 42.vecPK   ў,J�j�f�  W               �	 43.pPK   ў,J?P@s  �               � 43.vecPK   ў,J(���  [               w 44.pPK   ў,J���s  �               � 44.vecPK   ў,J�#�"  #               J 45.iPK   ў,J���  g               8 46.pPK   ў,J]��t  �               B< 46.vecPK   ў,J�Mx  �               �= 47.pPK   ў,J*s                 �A 47.vecPK   ў,J� �ӈ  �               BC 48.pPK   ў,J9u�u                 �F 48.vecPK   ў,J����  �               �H 49.pPK   ў,J�T�Os                 \L 49.vecPK   ў,J�%#�"  *#               N 50.iPK   ў,JG�M��  +               �p 51.pPK   ў,J[&��m                  �t 51.vecPK   ў,J�ғ�  \               jv 52.pPK   ў,J�;�s  �               �z 52.vecPK   ў,J��a  f               G| 53.pPK   ў,J���n  �               �� 53.vecPK   ў,J�}���  A               (� 54.pPK   ў,J�n��n  �               >� 54.vecPK   ў,J�gξ"  P#               �� 55.iPK   ў,J���                 Ъ 56.pPK   ў,J��3o                  �� 56.vecPK   ў,J�� �p  �               E� 57.pPK   ў,J���}p                 � 57.vecPK   ў,J�0���  5               �� 58.pPK   ў,J�1(Fp  �               �� 58.vecPK   ў,J�!��{  �               -� 59.pPK   ў,J�� �u                 ھ 59.vecPK   ў,J�[�#  �#               �� 60.iPK   ў,J��%�  :               �� 61.pPK   ў,JΞ�Cm                  �� 61.vecPK   ў,J�2��  @               u� 62.pPK   ў,J@w�4p                  �� 62.vecPK   ў,J���  >               (� 63.pPK   ў,J}Y��p                  7� 63.vecPK   ў,J*���  �               �� 64.pPK   ў,J9e�m                  �� 64.vecPK   ў,J5ר��"  Q#               F� 65.iPK   ў,J�T��  M               ; 66.pPK   ў,J�*`�m  �               ^! 66.vecPK   ў,J+�~�                 �" 67.pPK   ў,J�P]�q                  �& 67.vecPK   ў,JR2v  �               �( 68.pPK   ў,JNNRq                 *, 68.vecPK   ў,J�w��M  �               �- 69.pPK   ў,J���{w                 N1 69.vecPK   ў,Jv,_�"  7#               �2 70.iPK   ў,J�YQ�  �               �U 71.pPK   ў,Jԕ�"s                 �Y 71.vecPK   ў,J5�0]�  �               :[ 72.pPK   ў,J���\r                 �^ 72.vecPK   ў,J��^�  C               �` 73.pPK   ў,J��/1o                  �d 73.vecPK   ў,J���  ?               Df 74.pPK   ў,J,�q                  Zj 74.vecPK   ў,J�U0�"  9#               �k 75.iPK   ў,JED�o�  B               ܎ 76.pPK   ў,JSh�cn  �               � 76.vecPK   ў,J��H<�  I               �� 77.pPK   ў,J,Om  �               �� 77.vecPK   ў,JH�[>-  s               R� 78.pPK   ў,J���l  �               �� 78.vecPK   ў,Jӵ˰�                 Q� 79.pPK   ў,JY��'o                  6� 79.vecPK   ў,J���"  5#               ٥ 80.iPK   ў,J�@��                 �� 81.pPK   ў,J!�Ds                  �� 81.vecPK   ў,J��i�  9               >� 82.pPK   ў,J�+�>r  �               Y� 82.vecPK   ў,JC?�@�  A               �� 83.pPK   ў,J�2^p  �               � 83.vecPK   ў,J��  r               �� 84.pPK   ў,J@9�Bv  �               � 84.vecPK   ў,J5����"  �#               �� 85.iPK   ў,J	�2/  }               � 86.pPK   ў,Jj.�zs  �               @ 86.vecPK   ў,J��&/'  s               � 87.pPK   ў,J
��vu  �               @ 87.vecPK   ў,J
?�  _               � 88.pPK   ў,J���{s  �               ( 88.vecPK   ў,J��\�T  �               � 89.pPK   ў,J�N��n  �               U 89.vecPK   ў,J	�"  G#               � 90.iPK   ў,J���>�  I               �= 91.pPK   ў,JF#��s  �               B 91.vecPK   ў,J �_&�  A               �C 92.pPK   ў,JU�$by  �               �G 92.vecPK   ў,Jcyp��  9               yI 93.pPK   ў,J��u�q  �               �M 93.vecPK   ў,Jd�WU#  k               2O 94.pPK   ў,Js�r�r  �               �S 94.vecPK   ў,JYWE �"  �#               -U 95.iPK   ў,J��N�c  �               Tx 96.pPK   ў,J�T��m  �               �| 96.vecPK   ў,J��[k  �               �~ 97.pPK   ў,JSV6�l  �               '� 97.vecPK   ў,JT��)g  �               Ǆ 98.pPK   ў,Ju��n  �               `� 98.vecPK   ў,J\	���  �               � 99.pPK   ў,JFo�l  �               Ώ 99.vecPK   ў,JyF�Q#  �#               n� 100.iPK   ў,J����  �               �� 101.pPK   ў,J�2oxn  �               �� 101.vecPK   ў,JfۭV�  �               J� 102.pPK   ў,J�<'�p  �               � 102.vecPK   ў,J`�,  g               �� 103.pPK   ў,J7G�s  �               �� 103.vecPK   ў,J#k9(!  k               �� 104.pPK   ў,J`��km  �               �� 104.vecPK   ў,J��*�"  �#               �� 105.iPK   ў,Jl%Qb  �               �� 106.pPK   ў,J쨊�r  �               [� 106.vecPK   ў,J��1�  �               � 107.pPK   ў,J�X�k  �               �� 107.vecPK   ў,J�X�$�  �               o� 108.pPK   ў,JEB�%j  �               , 108.vecPK   ў,J�СF�  �               � 109.pPK   ў,JC�UXk  �               � 109.vecPK   ў,J#��#  �#               >
 110.iPK   ў,J����                 |- 111.pPK   ў,J��;um  �               v2 111.vecPK   ў,JV����  "               4 112.pPK   ў,J)z�h  �               ;9 112.vecPK   ў,J�����  �               �: 113.pPK   ў,J��Uch  �               �? 113.vecPK   ў,J�/�<�  �               nA 114.pPK   ў,J{�l  �               1F 114.vecPK   ў,J����"  b#               �G 115.iPK   ў,Jm;_T�  �               �j 116.pPK   ў,Jp�Jtm  �               �o 116.vecPK   ў,J<�]c�  �               4q 117.pPK   ў,J���j  �               5v 117.vecPK   ў,J>���  &               �w 118.pPK   ў,J���g  �               } 118.vecPK   ў,J�|�%  "               �~ 119.pPK   ў,JHJ�Uc  �               � 119.vecPK   ў,J>�M�"  $#               �� 120.iPK   ў,Jz�&�/  E               L� 121.pPK   ў,J,�<d  �               �� 121.vecPK   ў,J�Jt�  C               G� 122.pPK   ў,J�ǉtd  �               �� 122.vecPK   ў,Jy=u!r  �               -� 123.pPK   ў,J��b  �               һ 123.vecPK   ў,J{���  �               i� 124.pPK   ў,J���D^  �                � 124.vecPK   ў,J1 �t"   #               �� 125.iPK   ў,J�ݞ�                 Z� 126.pPK   ў,J_�<j  �               s� 126.vecPK   ў,J{+8�                 � 127.pPK   ў,J+Ҁ~h  �               !� 127.vecPK   ў,J猑��                 �� 128.pPK   ў,J�`��g  �               �� 128.vecPK   ў,J��A�;  N               v� 129.pPK   ў,J|n `  �               �  129.vecPK   ў,Jh�X"  �"               y 130.iPK   ў,J��#�*  >               % 131.pPK   ў,J��F�c  �               a* 131.vecPK   ў,Jǅ�u  3               �+ 132.pPK   ў,J��bUf  �               J1 132.vecPK   ў,J�Ê�e  p               �2 133.pPK   ў,J�pe�c  �               }8 133.vecPK   ў,J��K�m                 : 134.pPK   ў,J�FO^  �               �? 134.vecPK   ў,J�'/�2"  �"               HA 135.iPK   ў,J}�D��  �               �c 136.pPK   ў,J��FO\  �               �i 136.vecPK   ў,Jh��F~  �               k 137.pPK   ў,J#L+�b  �               �p 137.vecPK   ў,J��s�  *               \r 138.pPK   ў,J"��!o  �               �w 138.vecPK   ў,J�_?  /               @y 139.pPK   ў,Ju;6jl  �               �~ 139.vecPK   ў,J�r�!  ;"               *� 140.iPK   ў,J�yVi  s               	� 141.pPK   ў,J�vL�g  �               �� 141.vecPK   ў,J~���x  z               A� 142.pPK   ў,J�H�.c  �               � 142.vecPK   ў,JܧDY  a               �� 143.pPK   ў,J�k��i  �               � 143.vecPK   ў,J#ސ�  �               �� 144.pPK   ў,Jf��c  �               j� 144.vecPK   ў,J�+&�!  #"               � 145.iPK   ў,J��6i�  �               �� 146.pPK   ў,J�z`  �               �� 146.vecPK   ў,J'Y1��  �               V� 147.pPK   ў,J�eV�f  �               T� 147.vecPK   ў,J���  �               �� 148.pPK   ў,J�>��d  �               �� 148.vecPK   ў,J�X��  �               �� 149.pPK   ў,JJ�wUg  �               �� 149.vecPK   ў,Jxb��5!  �!               :� 150.iPK   ў,J{2Uщ  �               �  151.pPK   ў,J��ٙh  �               ^& 151.vecPK   ў,J���#�  �               �' 152.pPK   ў,J��Gc  �               �- 152.vecPK   ў,JJ��  �               �/ 153.pPK   ў,JS�0c  �               �5 153.vecPK   ў,J��p-�  �               I7 154.pPK   ў,J/��na  �               j= 154.vecPK   ў,J�/�B!  �!                ? 155.iPK   ў,J��#  	               u` 156.pPK   ў,J/;?b  �               �f 156.vecPK   ў,J�n��-  	               bh 157.pPK   ў,J\3��f  �               �n 157.vecPK   ў,Jq���  �               ]p 158.pPK   ў,Jy�kUa  �               �v 158.vecPK   ў,J��  �               <x 159.pPK   ў,J�kd  �               '~ 159.vecPK   ў,J�#�   �!               � 160.iPK   ў,J�0���  �               � 161.pPK   ў,J��f  �               � 161.vecPK   ў,J�+Փ�  �               �� 162.pPK   ў,J��-c  �               ۮ 162.vecPK   ў,JQ ��  �               s� 163.pPK   ў,J�a�k  �               �� 163.vecPK   ў,J
K�  �               ,� 164.pPK   ў,Jg&��g  �               0� 164.vecPK   ў,J/'!B�   J!               ̿ 165.iPK   ў,J�rC  ,	               �� 166.pPK   ў,JzXnd  �               0� 166.vecPK   ў,J�bծT  ;	               �� 167.pPK   ў,J�M*ed  �               P� 167.vecPK   ў,Jf䤅b  @	               �� 168.pPK   ў,JB�8*e  �               ~� 168.vecPK   ў,J:GF  +	               � 169.pPK   ў,J�b�Zc  �               �� 169.vecPK   ў,J�Y   �                ) 170.iPK   ў,J�KҬ  	               �! 171.pPK   ў,J/I2�j  �               �' 171.vecPK   ў,J��N�P  2	               �) 172.pPK   ў,J1AT�`  �               0 172.vecPK   ў,J�=�'^  =	               �1 173.pPK   ў,Jjm b  �               D8 173.vecPK   ў,J���  a	               �9 174.pPK   ў,Jk�9i  �               �@ 174.vecPK   ў,JnQ�   �                +B 175.iPK   ў,J֐�v4   	               kb 176.pPK   ў,J"q��g  �               �h 176.vecPK   ў,J��Ȓg  L	               nj 177.pPK   ў,J�#��g  �               q 177.vecPK   ў,J`a��  �	               �r 178.pPK   ў,J�Ia  �               �y 178.vecPK   ў,J�zMܺ  �	               { 179.pPK   ў,J�U��e  �               � 179.vecPK   ў,J�d�F�  d                �� 180.iPK   ў,Jdu��  m	               �� 181.pPK   ў,J�줔k  �               Z� 181.vecPK   ў,J�q?C�  e	               �� 182.pPK   ў,J>�ٲi  �               �� 182.vecPK   ў,J!;�`�  �	               M� 183.pPK   ў,JH�yd  �               =� 183.vecPK   ў,J��m�  �	               ּ 184.pPK   ў,J�3�c  �               �� 184.vecPK   ў,J�Wm  �               h� 185.iPK   ў,J�`��  �	               � 186.pPK   ў,J�Kd�f  �               � 186.vecPK   ў,Ji9� �  m	               �� 187.pPK   ў,JX}��k  �               r� 187.vecPK   ў,JD�ː�  n	               � 188.pPK   ў,J5�"�f  �               �� 188.vecPK   ў,JR	iu�  �	               q� 189.pPK   ў,J�O��d  �               s	 189.vecPK   ў,JGO:  �               	 190.iPK   ў,Jv�(�  �	               y&	 191.pPK   ў,JƗ��a  �               �-	 191.vecPK   ў,J����  �	               M/	 192.pPK   ў,J��v+e  �               [6	 192.vecPK   ў,J@b`�  �	               �7	 193.pPK   ў,J���d  �               �>	 193.vecPK   ў,J�p`U	  �	               �@	 194.pPK   ў,J��:�g  �               �G	 194.vecPK   ў,J���  �               gI	 195.iPK   ў,J���  �	               �h	 196.pPK   ў,J{:i`h  �               �o	 196.vecPK   ў,JFv�U  �	               pq	 197.pPK   ў,J�-�e  �               �x	 197.vecPK   ў,J��	�  �	               Xz	 198.pPK   ў,J�z8�h  �               ��	 198.vecPK   ў,J�5��  �	               :�	 199.pPK   ў,J�<,�e  �               k�	 199.vecPK   ў,J�W�}�  u               �	 200.iPK   ў,J�0�R  
               �	 201.pPK   ў,J�T�_`  �               ��	 201.vecPK   ў,JBeC�  R
               2�	 202.pPK   ў,J��ѡ^  �               �	 202.vecPK   ў,J�ߴ�S   
               ��	 203.pPK   ў,J#V�a  �               �	 203.vecPK   ў,JR�J�  F
               ��	 204.pPK   ў,J����`  �               `�	 204.vecPK   ў,J���  �               ��	 205.iPK   ў,JS�T�  �
               �	 206.pPK   ў,Ju�S�\  �               �	 206.vecPK   ў,J��� �  �
               ��	 207.pPK   ў,J�=(F`  �               � 
 207.vecPK   ў,J���  ^
               P
 208.pPK   ў,J���`  �               /

 208.vecPK   ў,J��ë�  Q
               �
 209.pPK   ў,Jruϓc  �               �
 209.vecPK   ў,J�zs�  <               )
 210.iPK   ў,J���  �
               4
 211.pPK   ў,J�:�b  �               <
 211.vecPK   ў,J}�X֢  ^
               �=
 212.pPK   ў,J�}8!b  �               zE
 212.vecPK   ў,J�0�  c
               G
 213.pPK   ў,J���d  �               �N
 213.vecPK   ў,J��c�  �
               wP
 214.pPK   ў,JpUE�a  �               �X
 214.vecPK   ў,J���<a  �               Z
 215.iPK   ў,J��Q�  m
               �x
 216.pPK   ў,J�IA�`  �               ��
 216.vecPK   ў,J���  �
               .�
 217.pPK   ў,JJ'��Y  �               G�
 217.vecPK   ў,JM֏�  �
               Ջ
 218.pPK   ў,J�q�m_  �               ד
 218.vecPK   ў,Jm�  �
               k�
 219.pPK   ў,J��n*\  �               ]�
 219.vecPK   ў,J�j��D  �               �
 220.iPK   ў,J�r3��  @
               e�
 221.pPK   ў,J��� ^  �               )�
 221.vecPK   ў,J�խ�}  2
               ��
 222.pPK   ў,JY�>�\  �               l�
 222.vecPK   ў,J�|i�  W
               ��
 223.pPK   ў,JI�K�_  �               ��
 223.vecPK   ў,J_��`�  n
               h�
 224.pPK   ў,J�l��^  �               Y�
 224.vecPK   ў,J�0�9�  P               ��
 225.iPK   ў,J\G�.�  �	               �  226.pPK   ў,J�YErj  �               � 226.vecPK   ў,J�K��  �	               �	 227.pPK   ў,J��@�e  �               � 227.vecPK   ў,J�*  �	               & 228.pPK   ў,J�"g  �               n 228.vecPK   ў,J$H  �	               
 229.pPK   ў,J׷%�h  �               N" 229.vecPK   ў,J���D  �               �# 230.iPK   ў,J���  �	               bA 231.pPK   ў,J��Nl  �               �H 231.vecPK   ў,J�'�*  �	               JJ 232.pPK   ў,Jg6�g  �               �Q 232.vecPK   ў,J���0  �	               S 233.pPK   ў,J8��c  �               �Z 233.vecPK   ў,JF7�h  '
               \ 234.pPK   ў,J�^�V[  �               �c 234.vecPK   ў,J��A��  �               Ee 235.iPK   ў,JQWu;  �	               r� 236.pPK   ў,J7��`  �               �� 236.vecPK   ў,JU7�q  ,
               u� 237.pPK   ў,J@T�9c  �               � 237.vecPK   ў,J\�J  
               �� 238.pPK   ў,J�2̺f  �               .� 238.vecPK   ў,J���C  

               ɝ 239.pPK   ў,Jt�m�h  �               ?� 239.vecPK    ��W  ܦ   